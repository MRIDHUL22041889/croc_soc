VERSION 5.7 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

PROPERTYDEFINITIONS
END PROPERTYDEFINITIONS


MACRO RM_IHPSG13_1P_256x64_c2_bm_bist
    CLASS BLOCK ;
    SIZE 784.48 BY 118.78 ;
    SYMMETRY X Y R90 ;
    PIN A_DIN[32]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  432.49 0 432.75 0.26 ;
        END
    END A_DIN[32]
    PIN A_DIN[31]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  351.73 0 351.99 0.26 ;
        END
    END A_DIN[31]
    PIN A_BIST_DIN[32]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  431.635 0 431.895 0.26 ;
        END
    END A_BIST_DIN[32]
    PIN A_BIST_DIN[31]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  352.585 0 352.845 0.26 ;
        END
    END A_BIST_DIN[31]
    PIN A_BM[32]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  424.65 0 424.91 0.26 ;
        END
    END A_BM[32]
    PIN A_BM[31]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  359.57 0 359.83 0.26 ;
        END
    END A_BM[31]
    PIN A_BIST_BM[32]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  426.025 0 426.285 0.26 ;
        END
    END A_BIST_BM[32]
    PIN A_BIST_BM[31]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  358.195 0 358.455 0.26 ;
        END
    END A_BIST_BM[31]
    PIN A_DOUT[32]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  425.16 0 425.42 0.26 ;
        END
    END A_DOUT[32]
    PIN A_DOUT[31]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  359.06 0 359.32 0.26 ;
        END
    END A_DOUT[31]
    PIN VSS!
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal4 ;
              RECT  771.79 0 774.6 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  760.55 0 763.36 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  749.31 0 752.12 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  738.07 0 740.88 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  726.83 0 729.64 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  715.59 0 718.4 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  704.35 0 707.16 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  693.11 0 695.92 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  681.87 0 684.68 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  670.63 0 673.44 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  659.39 0 662.2 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  648.15 0 650.96 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  636.91 0 639.72 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  625.67 0 628.48 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  614.43 0 617.24 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  603.19 0 606 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  591.95 0 594.76 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  580.71 0 583.52 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  569.47 0 572.28 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  558.23 0 561.04 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  546.99 0 549.8 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  535.75 0 538.56 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  524.51 0 527.32 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  513.27 0 516.08 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  502.03 0 504.84 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  490.79 0 493.6 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  479.55 0 482.36 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  468.31 0 471.12 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  457.07 0 459.88 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  445.83 0 448.64 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  434.59 0 437.4 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  423.35 0 426.16 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  408.86 0 411.67 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  398.56 0 401.37 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  383.11 0 385.92 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  372.81 0 375.62 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  358.32 0 361.13 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  347.08 0 349.89 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  335.84 0 338.65 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  324.6 0 327.41 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  313.36 0 316.17 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  302.12 0 304.93 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  290.88 0 293.69 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  279.64 0 282.45 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  268.4 0 271.21 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  257.16 0 259.97 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  245.92 0 248.73 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  234.68 0 237.49 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  223.44 0 226.25 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  212.2 0 215.01 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  200.96 0 203.77 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  189.72 0 192.53 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  178.48 0 181.29 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  167.24 0 170.05 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  156 0 158.81 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  144.76 0 147.57 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  133.52 0 136.33 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  122.28 0 125.09 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  111.04 0 113.85 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  99.8 0 102.61 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  88.56 0 91.37 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  77.32 0 80.13 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  66.08 0 68.89 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  54.84 0 57.65 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  43.6 0 46.41 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  32.36 0 35.17 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  21.12 0 23.93 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  9.88 0 12.69 118.78 ;
        END
    END VSS!
    PIN VDD!
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal4 ;
              RECT  777.41 0 780.22 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  766.17 0 768.98 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  754.93 0 757.74 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  743.69 0 746.5 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  732.45 0 735.26 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  721.21 0 724.02 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  709.97 0 712.78 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  698.73 0 701.54 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  687.49 0 690.3 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  676.25 0 679.06 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  665.01 0 667.82 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  653.77 0 656.58 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  642.53 0 645.34 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  631.29 0 634.1 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  620.05 0 622.86 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  608.81 0 611.62 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  597.57 0 600.38 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  586.33 0 589.14 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  575.09 0 577.9 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  563.85 0 566.66 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  552.61 0 555.42 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  541.37 0 544.18 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  530.13 0 532.94 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  518.89 0 521.7 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  507.65 0 510.46 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  496.41 0 499.22 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  485.17 0 487.98 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  473.93 0 476.74 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  462.69 0 465.5 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  451.45 0 454.26 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  440.21 0 443.02 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  428.97 0 431.78 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  403.71 0 406.52 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  393.41 0 396.22 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  388.26 0 391.07 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  377.96 0 380.77 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  352.7 0 355.51 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  341.46 0 344.27 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  330.22 0 333.03 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  318.98 0 321.79 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  307.74 0 310.55 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  296.5 0 299.31 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  285.26 0 288.07 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  274.02 0 276.83 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  262.78 0 265.59 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  251.54 0 254.35 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  240.3 0 243.11 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  229.06 0 231.87 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  217.82 0 220.63 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  206.58 0 209.39 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  195.34 0 198.15 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  184.1 0 186.91 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  172.86 0 175.67 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  161.62 0 164.43 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  150.38 0 153.19 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  139.14 0 141.95 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  127.9 0 130.71 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  116.66 0 119.47 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  105.42 0 108.23 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  94.18 0 96.99 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  82.94 0 85.75 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  71.7 0 74.51 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  60.46 0 63.27 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  49.22 0 52.03 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  37.98 0 40.79 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  26.74 0 29.55 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  15.5 0 18.31 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  4.26 0 7.07 38.825 ;
        END
    END VDD!
    PIN VDDARRAY!
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal4 ;
              RECT  777.41 45.465 780.22 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  766.17 45.465 768.98 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  754.93 45.465 757.74 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  743.69 45.465 746.5 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  732.45 45.465 735.26 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  721.21 45.465 724.02 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  709.97 45.465 712.78 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  698.73 45.465 701.54 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  687.49 45.465 690.3 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  676.25 45.465 679.06 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  665.01 45.465 667.82 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  653.77 45.465 656.58 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  642.53 45.465 645.34 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  631.29 45.465 634.1 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  620.05 45.465 622.86 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  608.81 45.465 611.62 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  597.57 45.465 600.38 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  586.33 45.465 589.14 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  575.09 45.465 577.9 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  563.85 45.465 566.66 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  552.61 45.465 555.42 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  541.37 45.465 544.18 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  530.13 45.465 532.94 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  518.89 45.465 521.7 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  507.65 45.465 510.46 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  496.41 45.465 499.22 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  485.17 45.465 487.98 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  473.93 45.465 476.74 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  462.69 45.465 465.5 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  451.45 45.465 454.26 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  440.21 45.465 443.02 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  428.97 45.465 431.78 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  352.7 45.465 355.51 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  341.46 45.465 344.27 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  330.22 45.465 333.03 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  318.98 45.465 321.79 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  307.74 45.465 310.55 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  296.5 45.465 299.31 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  285.26 45.465 288.07 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  274.02 45.465 276.83 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  262.78 45.465 265.59 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  251.54 45.465 254.35 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  240.3 45.465 243.11 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  229.06 45.465 231.87 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  217.82 45.465 220.63 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  206.58 45.465 209.39 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  195.34 45.465 198.15 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  184.1 45.465 186.91 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  172.86 45.465 175.67 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  161.62 45.465 164.43 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  150.38 45.465 153.19 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  139.14 45.465 141.95 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  127.9 45.465 130.71 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  116.66 45.465 119.47 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  105.42 45.465 108.23 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  94.18 45.465 96.99 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  82.94 45.465 85.75 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  71.7 45.465 74.51 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  60.46 45.465 63.27 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  49.22 45.465 52.03 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  37.98 45.465 40.79 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  26.74 45.465 29.55 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  15.5 45.465 18.31 118.78 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  4.26 45.465 7.07 118.78 ;
        END
    END VDDARRAY!
    PIN A_DIN[33]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  443.73 0 443.99 0.26 ;
        END
    END A_DIN[33]
    PIN A_DIN[30]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  340.49 0 340.75 0.26 ;
        END
    END A_DIN[30]
    PIN A_BIST_DIN[33]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  442.875 0 443.135 0.26 ;
        END
    END A_BIST_DIN[33]
    PIN A_BIST_DIN[30]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  341.345 0 341.605 0.26 ;
        END
    END A_BIST_DIN[30]
    PIN A_BM[33]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  435.89 0 436.15 0.26 ;
        END
    END A_BM[33]
    PIN A_BM[30]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  348.33 0 348.59 0.26 ;
        END
    END A_BM[30]
    PIN A_BIST_BM[33]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  437.265 0 437.525 0.26 ;
        END
    END A_BIST_BM[33]
    PIN A_BIST_BM[30]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  346.955 0 347.215 0.26 ;
        END
    END A_BIST_BM[30]
    PIN A_DOUT[33]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  436.4 0 436.66 0.26 ;
        END
    END A_DOUT[33]
    PIN A_DOUT[30]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  347.82 0 348.08 0.26 ;
        END
    END A_DOUT[30]
    PIN A_DIN[34]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  454.97 0 455.23 0.26 ;
        END
    END A_DIN[34]
    PIN A_DIN[29]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  329.25 0 329.51 0.26 ;
        END
    END A_DIN[29]
    PIN A_BIST_DIN[34]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  454.115 0 454.375 0.26 ;
        END
    END A_BIST_DIN[34]
    PIN A_BIST_DIN[29]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  330.105 0 330.365 0.26 ;
        END
    END A_BIST_DIN[29]
    PIN A_BM[34]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  447.13 0 447.39 0.26 ;
        END
    END A_BM[34]
    PIN A_BM[29]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  337.09 0 337.35 0.26 ;
        END
    END A_BM[29]
    PIN A_BIST_BM[34]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  448.505 0 448.765 0.26 ;
        END
    END A_BIST_BM[34]
    PIN A_BIST_BM[29]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  335.715 0 335.975 0.26 ;
        END
    END A_BIST_BM[29]
    PIN A_DOUT[34]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  447.64 0 447.9 0.26 ;
        END
    END A_DOUT[34]
    PIN A_DOUT[29]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  336.58 0 336.84 0.26 ;
        END
    END A_DOUT[29]
    PIN A_DIN[35]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  466.21 0 466.47 0.26 ;
        END
    END A_DIN[35]
    PIN A_DIN[28]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  318.01 0 318.27 0.26 ;
        END
    END A_DIN[28]
    PIN A_BIST_DIN[35]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  465.355 0 465.615 0.26 ;
        END
    END A_BIST_DIN[35]
    PIN A_BIST_DIN[28]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  318.865 0 319.125 0.26 ;
        END
    END A_BIST_DIN[28]
    PIN A_BM[35]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  458.37 0 458.63 0.26 ;
        END
    END A_BM[35]
    PIN A_BM[28]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  325.85 0 326.11 0.26 ;
        END
    END A_BM[28]
    PIN A_BIST_BM[35]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  459.745 0 460.005 0.26 ;
        END
    END A_BIST_BM[35]
    PIN A_BIST_BM[28]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  324.475 0 324.735 0.26 ;
        END
    END A_BIST_BM[28]
    PIN A_DOUT[35]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  458.88 0 459.14 0.26 ;
        END
    END A_DOUT[35]
    PIN A_DOUT[28]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  325.34 0 325.6 0.26 ;
        END
    END A_DOUT[28]
    PIN A_DIN[36]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  477.45 0 477.71 0.26 ;
        END
    END A_DIN[36]
    PIN A_DIN[27]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  306.77 0 307.03 0.26 ;
        END
    END A_DIN[27]
    PIN A_BIST_DIN[36]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  476.595 0 476.855 0.26 ;
        END
    END A_BIST_DIN[36]
    PIN A_BIST_DIN[27]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  307.625 0 307.885 0.26 ;
        END
    END A_BIST_DIN[27]
    PIN A_BM[36]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  469.61 0 469.87 0.26 ;
        END
    END A_BM[36]
    PIN A_BM[27]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  314.61 0 314.87 0.26 ;
        END
    END A_BM[27]
    PIN A_BIST_BM[36]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  470.985 0 471.245 0.26 ;
        END
    END A_BIST_BM[36]
    PIN A_BIST_BM[27]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  313.235 0 313.495 0.26 ;
        END
    END A_BIST_BM[27]
    PIN A_DOUT[36]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  470.12 0 470.38 0.26 ;
        END
    END A_DOUT[36]
    PIN A_DOUT[27]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  314.1 0 314.36 0.26 ;
        END
    END A_DOUT[27]
    PIN A_DIN[37]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  488.69 0 488.95 0.26 ;
        END
    END A_DIN[37]
    PIN A_DIN[26]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  295.53 0 295.79 0.26 ;
        END
    END A_DIN[26]
    PIN A_BIST_DIN[37]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  487.835 0 488.095 0.26 ;
        END
    END A_BIST_DIN[37]
    PIN A_BIST_DIN[26]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  296.385 0 296.645 0.26 ;
        END
    END A_BIST_DIN[26]
    PIN A_BM[37]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  480.85 0 481.11 0.26 ;
        END
    END A_BM[37]
    PIN A_BM[26]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  303.37 0 303.63 0.26 ;
        END
    END A_BM[26]
    PIN A_BIST_BM[37]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  482.225 0 482.485 0.26 ;
        END
    END A_BIST_BM[37]
    PIN A_BIST_BM[26]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  301.995 0 302.255 0.26 ;
        END
    END A_BIST_BM[26]
    PIN A_DOUT[37]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  481.36 0 481.62 0.26 ;
        END
    END A_DOUT[37]
    PIN A_DOUT[26]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  302.86 0 303.12 0.26 ;
        END
    END A_DOUT[26]
    PIN A_DIN[38]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  499.93 0 500.19 0.26 ;
        END
    END A_DIN[38]
    PIN A_DIN[25]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  284.29 0 284.55 0.26 ;
        END
    END A_DIN[25]
    PIN A_BIST_DIN[38]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  499.075 0 499.335 0.26 ;
        END
    END A_BIST_DIN[38]
    PIN A_BIST_DIN[25]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  285.145 0 285.405 0.26 ;
        END
    END A_BIST_DIN[25]
    PIN A_BM[38]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  492.09 0 492.35 0.26 ;
        END
    END A_BM[38]
    PIN A_BM[25]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  292.13 0 292.39 0.26 ;
        END
    END A_BM[25]
    PIN A_BIST_BM[38]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  493.465 0 493.725 0.26 ;
        END
    END A_BIST_BM[38]
    PIN A_BIST_BM[25]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  290.755 0 291.015 0.26 ;
        END
    END A_BIST_BM[25]
    PIN A_DOUT[38]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  492.6 0 492.86 0.26 ;
        END
    END A_DOUT[38]
    PIN A_DOUT[25]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  291.62 0 291.88 0.26 ;
        END
    END A_DOUT[25]
    PIN A_DIN[39]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  511.17 0 511.43 0.26 ;
        END
    END A_DIN[39]
    PIN A_DIN[24]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  273.05 0 273.31 0.26 ;
        END
    END A_DIN[24]
    PIN A_BIST_DIN[39]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  510.315 0 510.575 0.26 ;
        END
    END A_BIST_DIN[39]
    PIN A_BIST_DIN[24]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  273.905 0 274.165 0.26 ;
        END
    END A_BIST_DIN[24]
    PIN A_BM[39]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  503.33 0 503.59 0.26 ;
        END
    END A_BM[39]
    PIN A_BM[24]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  280.89 0 281.15 0.26 ;
        END
    END A_BM[24]
    PIN A_BIST_BM[39]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  504.705 0 504.965 0.26 ;
        END
    END A_BIST_BM[39]
    PIN A_BIST_BM[24]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  279.515 0 279.775 0.26 ;
        END
    END A_BIST_BM[24]
    PIN A_DOUT[39]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  503.84 0 504.1 0.26 ;
        END
    END A_DOUT[39]
    PIN A_DOUT[24]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  280.38 0 280.64 0.26 ;
        END
    END A_DOUT[24]
    PIN A_DIN[40]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  522.41 0 522.67 0.26 ;
        END
    END A_DIN[40]
    PIN A_DIN[23]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  261.81 0 262.07 0.26 ;
        END
    END A_DIN[23]
    PIN A_BIST_DIN[40]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  521.555 0 521.815 0.26 ;
        END
    END A_BIST_DIN[40]
    PIN A_BIST_DIN[23]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  262.665 0 262.925 0.26 ;
        END
    END A_BIST_DIN[23]
    PIN A_BM[40]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  514.57 0 514.83 0.26 ;
        END
    END A_BM[40]
    PIN A_BM[23]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  269.65 0 269.91 0.26 ;
        END
    END A_BM[23]
    PIN A_BIST_BM[40]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  515.945 0 516.205 0.26 ;
        END
    END A_BIST_BM[40]
    PIN A_BIST_BM[23]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  268.275 0 268.535 0.26 ;
        END
    END A_BIST_BM[23]
    PIN A_DOUT[40]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  515.08 0 515.34 0.26 ;
        END
    END A_DOUT[40]
    PIN A_DOUT[23]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  269.14 0 269.4 0.26 ;
        END
    END A_DOUT[23]
    PIN A_DIN[41]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  533.65 0 533.91 0.26 ;
        END
    END A_DIN[41]
    PIN A_DIN[22]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  250.57 0 250.83 0.26 ;
        END
    END A_DIN[22]
    PIN A_BIST_DIN[41]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  532.795 0 533.055 0.26 ;
        END
    END A_BIST_DIN[41]
    PIN A_BIST_DIN[22]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  251.425 0 251.685 0.26 ;
        END
    END A_BIST_DIN[22]
    PIN A_BM[41]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  525.81 0 526.07 0.26 ;
        END
    END A_BM[41]
    PIN A_BM[22]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  258.41 0 258.67 0.26 ;
        END
    END A_BM[22]
    PIN A_BIST_BM[41]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  527.185 0 527.445 0.26 ;
        END
    END A_BIST_BM[41]
    PIN A_BIST_BM[22]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  257.035 0 257.295 0.26 ;
        END
    END A_BIST_BM[22]
    PIN A_DOUT[41]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  526.32 0 526.58 0.26 ;
        END
    END A_DOUT[41]
    PIN A_DOUT[22]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  257.9 0 258.16 0.26 ;
        END
    END A_DOUT[22]
    PIN A_DIN[42]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  544.89 0 545.15 0.26 ;
        END
    END A_DIN[42]
    PIN A_DIN[21]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  239.33 0 239.59 0.26 ;
        END
    END A_DIN[21]
    PIN A_BIST_DIN[42]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  544.035 0 544.295 0.26 ;
        END
    END A_BIST_DIN[42]
    PIN A_BIST_DIN[21]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  240.185 0 240.445 0.26 ;
        END
    END A_BIST_DIN[21]
    PIN A_BM[42]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  537.05 0 537.31 0.26 ;
        END
    END A_BM[42]
    PIN A_BM[21]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  247.17 0 247.43 0.26 ;
        END
    END A_BM[21]
    PIN A_BIST_BM[42]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  538.425 0 538.685 0.26 ;
        END
    END A_BIST_BM[42]
    PIN A_BIST_BM[21]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  245.795 0 246.055 0.26 ;
        END
    END A_BIST_BM[21]
    PIN A_DOUT[42]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  537.56 0 537.82 0.26 ;
        END
    END A_DOUT[42]
    PIN A_DOUT[21]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  246.66 0 246.92 0.26 ;
        END
    END A_DOUT[21]
    PIN A_DIN[43]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  556.13 0 556.39 0.26 ;
        END
    END A_DIN[43]
    PIN A_DIN[20]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  228.09 0 228.35 0.26 ;
        END
    END A_DIN[20]
    PIN A_BIST_DIN[43]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  555.275 0 555.535 0.26 ;
        END
    END A_BIST_DIN[43]
    PIN A_BIST_DIN[20]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  228.945 0 229.205 0.26 ;
        END
    END A_BIST_DIN[20]
    PIN A_BM[43]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  548.29 0 548.55 0.26 ;
        END
    END A_BM[43]
    PIN A_BM[20]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  235.93 0 236.19 0.26 ;
        END
    END A_BM[20]
    PIN A_BIST_BM[43]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  549.665 0 549.925 0.26 ;
        END
    END A_BIST_BM[43]
    PIN A_BIST_BM[20]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  234.555 0 234.815 0.26 ;
        END
    END A_BIST_BM[20]
    PIN A_DOUT[43]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  548.8 0 549.06 0.26 ;
        END
    END A_DOUT[43]
    PIN A_DOUT[20]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  235.42 0 235.68 0.26 ;
        END
    END A_DOUT[20]
    PIN A_DIN[44]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  567.37 0 567.63 0.26 ;
        END
    END A_DIN[44]
    PIN A_DIN[19]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  216.85 0 217.11 0.26 ;
        END
    END A_DIN[19]
    PIN A_BIST_DIN[44]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  566.515 0 566.775 0.26 ;
        END
    END A_BIST_DIN[44]
    PIN A_BIST_DIN[19]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  217.705 0 217.965 0.26 ;
        END
    END A_BIST_DIN[19]
    PIN A_BM[44]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  559.53 0 559.79 0.26 ;
        END
    END A_BM[44]
    PIN A_BM[19]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  224.69 0 224.95 0.26 ;
        END
    END A_BM[19]
    PIN A_BIST_BM[44]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  560.905 0 561.165 0.26 ;
        END
    END A_BIST_BM[44]
    PIN A_BIST_BM[19]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  223.315 0 223.575 0.26 ;
        END
    END A_BIST_BM[19]
    PIN A_DOUT[44]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  560.04 0 560.3 0.26 ;
        END
    END A_DOUT[44]
    PIN A_DOUT[19]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  224.18 0 224.44 0.26 ;
        END
    END A_DOUT[19]
    PIN A_DIN[45]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  578.61 0 578.87 0.26 ;
        END
    END A_DIN[45]
    PIN A_DIN[18]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  205.61 0 205.87 0.26 ;
        END
    END A_DIN[18]
    PIN A_BIST_DIN[45]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  577.755 0 578.015 0.26 ;
        END
    END A_BIST_DIN[45]
    PIN A_BIST_DIN[18]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  206.465 0 206.725 0.26 ;
        END
    END A_BIST_DIN[18]
    PIN A_BM[45]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  570.77 0 571.03 0.26 ;
        END
    END A_BM[45]
    PIN A_BM[18]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  213.45 0 213.71 0.26 ;
        END
    END A_BM[18]
    PIN A_BIST_BM[45]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  572.145 0 572.405 0.26 ;
        END
    END A_BIST_BM[45]
    PIN A_BIST_BM[18]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  212.075 0 212.335 0.26 ;
        END
    END A_BIST_BM[18]
    PIN A_DOUT[45]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  571.28 0 571.54 0.26 ;
        END
    END A_DOUT[45]
    PIN A_DOUT[18]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  212.94 0 213.2 0.26 ;
        END
    END A_DOUT[18]
    PIN A_DIN[46]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  589.85 0 590.11 0.26 ;
        END
    END A_DIN[46]
    PIN A_DIN[17]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  194.37 0 194.63 0.26 ;
        END
    END A_DIN[17]
    PIN A_BIST_DIN[46]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  588.995 0 589.255 0.26 ;
        END
    END A_BIST_DIN[46]
    PIN A_BIST_DIN[17]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  195.225 0 195.485 0.26 ;
        END
    END A_BIST_DIN[17]
    PIN A_BM[46]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  582.01 0 582.27 0.26 ;
        END
    END A_BM[46]
    PIN A_BM[17]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  202.21 0 202.47 0.26 ;
        END
    END A_BM[17]
    PIN A_BIST_BM[46]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  583.385 0 583.645 0.26 ;
        END
    END A_BIST_BM[46]
    PIN A_BIST_BM[17]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  200.835 0 201.095 0.26 ;
        END
    END A_BIST_BM[17]
    PIN A_DOUT[46]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  582.52 0 582.78 0.26 ;
        END
    END A_DOUT[46]
    PIN A_DOUT[17]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  201.7 0 201.96 0.26 ;
        END
    END A_DOUT[17]
    PIN A_DIN[47]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  601.09 0 601.35 0.26 ;
        END
    END A_DIN[47]
    PIN A_DIN[16]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  183.13 0 183.39 0.26 ;
        END
    END A_DIN[16]
    PIN A_BIST_DIN[47]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  600.235 0 600.495 0.26 ;
        END
    END A_BIST_DIN[47]
    PIN A_BIST_DIN[16]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  183.985 0 184.245 0.26 ;
        END
    END A_BIST_DIN[16]
    PIN A_BM[47]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  593.25 0 593.51 0.26 ;
        END
    END A_BM[47]
    PIN A_BM[16]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  190.97 0 191.23 0.26 ;
        END
    END A_BM[16]
    PIN A_BIST_BM[47]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  594.625 0 594.885 0.26 ;
        END
    END A_BIST_BM[47]
    PIN A_BIST_BM[16]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  189.595 0 189.855 0.26 ;
        END
    END A_BIST_BM[16]
    PIN A_DOUT[47]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  593.76 0 594.02 0.26 ;
        END
    END A_DOUT[47]
    PIN A_DOUT[16]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  190.46 0 190.72 0.26 ;
        END
    END A_DOUT[16]
    PIN A_DIN[48]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  612.33 0 612.59 0.26 ;
        END
    END A_DIN[48]
    PIN A_DIN[15]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  171.89 0 172.15 0.26 ;
        END
    END A_DIN[15]
    PIN A_BIST_DIN[48]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  611.475 0 611.735 0.26 ;
        END
    END A_BIST_DIN[48]
    PIN A_BIST_DIN[15]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  172.745 0 173.005 0.26 ;
        END
    END A_BIST_DIN[15]
    PIN A_BM[48]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  604.49 0 604.75 0.26 ;
        END
    END A_BM[48]
    PIN A_BM[15]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  179.73 0 179.99 0.26 ;
        END
    END A_BM[15]
    PIN A_BIST_BM[48]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  605.865 0 606.125 0.26 ;
        END
    END A_BIST_BM[48]
    PIN A_BIST_BM[15]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  178.355 0 178.615 0.26 ;
        END
    END A_BIST_BM[15]
    PIN A_DOUT[48]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  605 0 605.26 0.26 ;
        END
    END A_DOUT[48]
    PIN A_DOUT[15]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  179.22 0 179.48 0.26 ;
        END
    END A_DOUT[15]
    PIN A_DIN[49]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  623.57 0 623.83 0.26 ;
        END
    END A_DIN[49]
    PIN A_DIN[14]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  160.65 0 160.91 0.26 ;
        END
    END A_DIN[14]
    PIN A_BIST_DIN[49]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  622.715 0 622.975 0.26 ;
        END
    END A_BIST_DIN[49]
    PIN A_BIST_DIN[14]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  161.505 0 161.765 0.26 ;
        END
    END A_BIST_DIN[14]
    PIN A_BM[49]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  615.73 0 615.99 0.26 ;
        END
    END A_BM[49]
    PIN A_BM[14]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  168.49 0 168.75 0.26 ;
        END
    END A_BM[14]
    PIN A_BIST_BM[49]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  617.105 0 617.365 0.26 ;
        END
    END A_BIST_BM[49]
    PIN A_BIST_BM[14]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  167.115 0 167.375 0.26 ;
        END
    END A_BIST_BM[14]
    PIN A_DOUT[49]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  616.24 0 616.5 0.26 ;
        END
    END A_DOUT[49]
    PIN A_DOUT[14]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  167.98 0 168.24 0.26 ;
        END
    END A_DOUT[14]
    PIN A_DIN[50]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  634.81 0 635.07 0.26 ;
        END
    END A_DIN[50]
    PIN A_DIN[13]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  149.41 0 149.67 0.26 ;
        END
    END A_DIN[13]
    PIN A_BIST_DIN[50]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  633.955 0 634.215 0.26 ;
        END
    END A_BIST_DIN[50]
    PIN A_BIST_DIN[13]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  150.265 0 150.525 0.26 ;
        END
    END A_BIST_DIN[13]
    PIN A_BM[50]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  626.97 0 627.23 0.26 ;
        END
    END A_BM[50]
    PIN A_BM[13]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  157.25 0 157.51 0.26 ;
        END
    END A_BM[13]
    PIN A_BIST_BM[50]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  628.345 0 628.605 0.26 ;
        END
    END A_BIST_BM[50]
    PIN A_BIST_BM[13]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  155.875 0 156.135 0.26 ;
        END
    END A_BIST_BM[13]
    PIN A_DOUT[50]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  627.48 0 627.74 0.26 ;
        END
    END A_DOUT[50]
    PIN A_DOUT[13]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  156.74 0 157 0.26 ;
        END
    END A_DOUT[13]
    PIN A_DIN[51]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  646.05 0 646.31 0.26 ;
        END
    END A_DIN[51]
    PIN A_DIN[12]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  138.17 0 138.43 0.26 ;
        END
    END A_DIN[12]
    PIN A_BIST_DIN[51]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  645.195 0 645.455 0.26 ;
        END
    END A_BIST_DIN[51]
    PIN A_BIST_DIN[12]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  139.025 0 139.285 0.26 ;
        END
    END A_BIST_DIN[12]
    PIN A_BM[51]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  638.21 0 638.47 0.26 ;
        END
    END A_BM[51]
    PIN A_BM[12]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  146.01 0 146.27 0.26 ;
        END
    END A_BM[12]
    PIN A_BIST_BM[51]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  639.585 0 639.845 0.26 ;
        END
    END A_BIST_BM[51]
    PIN A_BIST_BM[12]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  144.635 0 144.895 0.26 ;
        END
    END A_BIST_BM[12]
    PIN A_DOUT[51]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  638.72 0 638.98 0.26 ;
        END
    END A_DOUT[51]
    PIN A_DOUT[12]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  145.5 0 145.76 0.26 ;
        END
    END A_DOUT[12]
    PIN A_DIN[52]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  657.29 0 657.55 0.26 ;
        END
    END A_DIN[52]
    PIN A_DIN[11]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  126.93 0 127.19 0.26 ;
        END
    END A_DIN[11]
    PIN A_BIST_DIN[52]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  656.435 0 656.695 0.26 ;
        END
    END A_BIST_DIN[52]
    PIN A_BIST_DIN[11]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  127.785 0 128.045 0.26 ;
        END
    END A_BIST_DIN[11]
    PIN A_BM[52]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  649.45 0 649.71 0.26 ;
        END
    END A_BM[52]
    PIN A_BM[11]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  134.77 0 135.03 0.26 ;
        END
    END A_BM[11]
    PIN A_BIST_BM[52]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  650.825 0 651.085 0.26 ;
        END
    END A_BIST_BM[52]
    PIN A_BIST_BM[11]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  133.395 0 133.655 0.26 ;
        END
    END A_BIST_BM[11]
    PIN A_DOUT[52]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  649.96 0 650.22 0.26 ;
        END
    END A_DOUT[52]
    PIN A_DOUT[11]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  134.26 0 134.52 0.26 ;
        END
    END A_DOUT[11]
    PIN A_DIN[53]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  668.53 0 668.79 0.26 ;
        END
    END A_DIN[53]
    PIN A_DIN[10]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  115.69 0 115.95 0.26 ;
        END
    END A_DIN[10]
    PIN A_BIST_DIN[53]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  667.675 0 667.935 0.26 ;
        END
    END A_BIST_DIN[53]
    PIN A_BIST_DIN[10]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  116.545 0 116.805 0.26 ;
        END
    END A_BIST_DIN[10]
    PIN A_BM[53]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  660.69 0 660.95 0.26 ;
        END
    END A_BM[53]
    PIN A_BM[10]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  123.53 0 123.79 0.26 ;
        END
    END A_BM[10]
    PIN A_BIST_BM[53]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  662.065 0 662.325 0.26 ;
        END
    END A_BIST_BM[53]
    PIN A_BIST_BM[10]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  122.155 0 122.415 0.26 ;
        END
    END A_BIST_BM[10]
    PIN A_DOUT[53]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  661.2 0 661.46 0.26 ;
        END
    END A_DOUT[53]
    PIN A_DOUT[10]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  123.02 0 123.28 0.26 ;
        END
    END A_DOUT[10]
    PIN A_DIN[54]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  679.77 0 680.03 0.26 ;
        END
    END A_DIN[54]
    PIN A_DIN[9]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  104.45 0 104.71 0.26 ;
        END
    END A_DIN[9]
    PIN A_BIST_DIN[54]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  678.915 0 679.175 0.26 ;
        END
    END A_BIST_DIN[54]
    PIN A_BIST_DIN[9]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  105.305 0 105.565 0.26 ;
        END
    END A_BIST_DIN[9]
    PIN A_BM[54]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  671.93 0 672.19 0.26 ;
        END
    END A_BM[54]
    PIN A_BM[9]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  112.29 0 112.55 0.26 ;
        END
    END A_BM[9]
    PIN A_BIST_BM[54]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  673.305 0 673.565 0.26 ;
        END
    END A_BIST_BM[54]
    PIN A_BIST_BM[9]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  110.915 0 111.175 0.26 ;
        END
    END A_BIST_BM[9]
    PIN A_DOUT[54]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  672.44 0 672.7 0.26 ;
        END
    END A_DOUT[54]
    PIN A_DOUT[9]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  111.78 0 112.04 0.26 ;
        END
    END A_DOUT[9]
    PIN A_DIN[55]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  691.01 0 691.27 0.26 ;
        END
    END A_DIN[55]
    PIN A_DIN[8]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  93.21 0 93.47 0.26 ;
        END
    END A_DIN[8]
    PIN A_BIST_DIN[55]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  690.155 0 690.415 0.26 ;
        END
    END A_BIST_DIN[55]
    PIN A_BIST_DIN[8]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  94.065 0 94.325 0.26 ;
        END
    END A_BIST_DIN[8]
    PIN A_BM[55]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  683.17 0 683.43 0.26 ;
        END
    END A_BM[55]
    PIN A_BM[8]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  101.05 0 101.31 0.26 ;
        END
    END A_BM[8]
    PIN A_BIST_BM[55]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  684.545 0 684.805 0.26 ;
        END
    END A_BIST_BM[55]
    PIN A_BIST_BM[8]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  99.675 0 99.935 0.26 ;
        END
    END A_BIST_BM[8]
    PIN A_DOUT[55]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  683.68 0 683.94 0.26 ;
        END
    END A_DOUT[55]
    PIN A_DOUT[8]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  100.54 0 100.8 0.26 ;
        END
    END A_DOUT[8]
    PIN A_DIN[56]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  702.25 0 702.51 0.26 ;
        END
    END A_DIN[56]
    PIN A_DIN[7]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  81.97 0 82.23 0.26 ;
        END
    END A_DIN[7]
    PIN A_BIST_DIN[56]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  701.395 0 701.655 0.26 ;
        END
    END A_BIST_DIN[56]
    PIN A_BIST_DIN[7]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  82.825 0 83.085 0.26 ;
        END
    END A_BIST_DIN[7]
    PIN A_BM[56]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  694.41 0 694.67 0.26 ;
        END
    END A_BM[56]
    PIN A_BM[7]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  89.81 0 90.07 0.26 ;
        END
    END A_BM[7]
    PIN A_BIST_BM[56]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  695.785 0 696.045 0.26 ;
        END
    END A_BIST_BM[56]
    PIN A_BIST_BM[7]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  88.435 0 88.695 0.26 ;
        END
    END A_BIST_BM[7]
    PIN A_DOUT[56]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  694.92 0 695.18 0.26 ;
        END
    END A_DOUT[56]
    PIN A_DOUT[7]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  89.3 0 89.56 0.26 ;
        END
    END A_DOUT[7]
    PIN A_DIN[57]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  713.49 0 713.75 0.26 ;
        END
    END A_DIN[57]
    PIN A_DIN[6]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  70.73 0 70.99 0.26 ;
        END
    END A_DIN[6]
    PIN A_BIST_DIN[57]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  712.635 0 712.895 0.26 ;
        END
    END A_BIST_DIN[57]
    PIN A_BIST_DIN[6]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  71.585 0 71.845 0.26 ;
        END
    END A_BIST_DIN[6]
    PIN A_BM[57]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  705.65 0 705.91 0.26 ;
        END
    END A_BM[57]
    PIN A_BM[6]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  78.57 0 78.83 0.26 ;
        END
    END A_BM[6]
    PIN A_BIST_BM[57]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  707.025 0 707.285 0.26 ;
        END
    END A_BIST_BM[57]
    PIN A_BIST_BM[6]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  77.195 0 77.455 0.26 ;
        END
    END A_BIST_BM[6]
    PIN A_DOUT[57]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  706.16 0 706.42 0.26 ;
        END
    END A_DOUT[57]
    PIN A_DOUT[6]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  78.06 0 78.32 0.26 ;
        END
    END A_DOUT[6]
    PIN A_DIN[58]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  724.73 0 724.99 0.26 ;
        END
    END A_DIN[58]
    PIN A_DIN[5]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  59.49 0 59.75 0.26 ;
        END
    END A_DIN[5]
    PIN A_BIST_DIN[58]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  723.875 0 724.135 0.26 ;
        END
    END A_BIST_DIN[58]
    PIN A_BIST_DIN[5]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  60.345 0 60.605 0.26 ;
        END
    END A_BIST_DIN[5]
    PIN A_BM[58]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  716.89 0 717.15 0.26 ;
        END
    END A_BM[58]
    PIN A_BM[5]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  67.33 0 67.59 0.26 ;
        END
    END A_BM[5]
    PIN A_BIST_BM[58]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  718.265 0 718.525 0.26 ;
        END
    END A_BIST_BM[58]
    PIN A_BIST_BM[5]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  65.955 0 66.215 0.26 ;
        END
    END A_BIST_BM[5]
    PIN A_DOUT[58]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  717.4 0 717.66 0.26 ;
        END
    END A_DOUT[58]
    PIN A_DOUT[5]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  66.82 0 67.08 0.26 ;
        END
    END A_DOUT[5]
    PIN A_DIN[59]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  735.97 0 736.23 0.26 ;
        END
    END A_DIN[59]
    PIN A_DIN[4]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  48.25 0 48.51 0.26 ;
        END
    END A_DIN[4]
    PIN A_BIST_DIN[59]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  735.115 0 735.375 0.26 ;
        END
    END A_BIST_DIN[59]
    PIN A_BIST_DIN[4]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  49.105 0 49.365 0.26 ;
        END
    END A_BIST_DIN[4]
    PIN A_BM[59]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  728.13 0 728.39 0.26 ;
        END
    END A_BM[59]
    PIN A_BM[4]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  56.09 0 56.35 0.26 ;
        END
    END A_BM[4]
    PIN A_BIST_BM[59]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  729.505 0 729.765 0.26 ;
        END
    END A_BIST_BM[59]
    PIN A_BIST_BM[4]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  54.715 0 54.975 0.26 ;
        END
    END A_BIST_BM[4]
    PIN A_DOUT[59]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  728.64 0 728.9 0.26 ;
        END
    END A_DOUT[59]
    PIN A_DOUT[4]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  55.58 0 55.84 0.26 ;
        END
    END A_DOUT[4]
    PIN A_DIN[60]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  747.21 0 747.47 0.26 ;
        END
    END A_DIN[60]
    PIN A_DIN[3]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  37.01 0 37.27 0.26 ;
        END
    END A_DIN[3]
    PIN A_BIST_DIN[60]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  746.355 0 746.615 0.26 ;
        END
    END A_BIST_DIN[60]
    PIN A_BIST_DIN[3]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  37.865 0 38.125 0.26 ;
        END
    END A_BIST_DIN[3]
    PIN A_BM[60]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  739.37 0 739.63 0.26 ;
        END
    END A_BM[60]
    PIN A_BM[3]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  44.85 0 45.11 0.26 ;
        END
    END A_BM[3]
    PIN A_BIST_BM[60]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  740.745 0 741.005 0.26 ;
        END
    END A_BIST_BM[60]
    PIN A_BIST_BM[3]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  43.475 0 43.735 0.26 ;
        END
    END A_BIST_BM[3]
    PIN A_DOUT[60]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  739.88 0 740.14 0.26 ;
        END
    END A_DOUT[60]
    PIN A_DOUT[3]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  44.34 0 44.6 0.26 ;
        END
    END A_DOUT[3]
    PIN A_DIN[61]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  758.45 0 758.71 0.26 ;
        END
    END A_DIN[61]
    PIN A_DIN[2]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  25.77 0 26.03 0.26 ;
        END
    END A_DIN[2]
    PIN A_BIST_DIN[61]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  757.595 0 757.855 0.26 ;
        END
    END A_BIST_DIN[61]
    PIN A_BIST_DIN[2]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  26.625 0 26.885 0.26 ;
        END
    END A_BIST_DIN[2]
    PIN A_BM[61]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  750.61 0 750.87 0.26 ;
        END
    END A_BM[61]
    PIN A_BM[2]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  33.61 0 33.87 0.26 ;
        END
    END A_BM[2]
    PIN A_BIST_BM[61]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  751.985 0 752.245 0.26 ;
        END
    END A_BIST_BM[61]
    PIN A_BIST_BM[2]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  32.235 0 32.495 0.26 ;
        END
    END A_BIST_BM[2]
    PIN A_DOUT[61]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  751.12 0 751.38 0.26 ;
        END
    END A_DOUT[61]
    PIN A_DOUT[2]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  33.1 0 33.36 0.26 ;
        END
    END A_DOUT[2]
    PIN A_DIN[62]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  769.69 0 769.95 0.26 ;
        END
    END A_DIN[62]
    PIN A_DIN[1]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  14.53 0 14.79 0.26 ;
        END
    END A_DIN[1]
    PIN A_BIST_DIN[62]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  768.835 0 769.095 0.26 ;
        END
    END A_BIST_DIN[62]
    PIN A_BIST_DIN[1]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  15.385 0 15.645 0.26 ;
        END
    END A_BIST_DIN[1]
    PIN A_BM[62]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  761.85 0 762.11 0.26 ;
        END
    END A_BM[62]
    PIN A_BM[1]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  22.37 0 22.63 0.26 ;
        END
    END A_BM[1]
    PIN A_BIST_BM[62]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  763.225 0 763.485 0.26 ;
        END
    END A_BIST_BM[62]
    PIN A_BIST_BM[1]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  20.995 0 21.255 0.26 ;
        END
    END A_BIST_BM[1]
    PIN A_DOUT[62]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  762.36 0 762.62 0.26 ;
        END
    END A_DOUT[62]
    PIN A_DOUT[1]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  21.86 0 22.12 0.26 ;
        END
    END A_DOUT[1]
    PIN A_DIN[63]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  780.93 0 781.19 0.26 ;
        END
    END A_DIN[63]
    PIN A_DIN[0]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  3.29 0 3.55 0.26 ;
        END
    END A_DIN[0]
    PIN A_BIST_DIN[63]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  780.075 0 780.335 0.26 ;
        END
    END A_BIST_DIN[63]
    PIN A_BIST_DIN[0]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  4.145 0 4.405 0.26 ;
        END
    END A_BIST_DIN[0]
    PIN A_BM[63]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  773.09 0 773.35 0.26 ;
        END
    END A_BM[63]
    PIN A_BM[0]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  11.13 0 11.39 0.26 ;
        END
    END A_BM[0]
    PIN A_BIST_BM[63]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  774.465 0 774.725 0.26 ;
        END
    END A_BIST_BM[63]
    PIN A_BIST_BM[0]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  9.755 0 10.015 0.26 ;
        END
    END A_BIST_BM[0]
    PIN A_DOUT[63]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  773.6 0 773.86 0.26 ;
        END
    END A_DOUT[63]
    PIN A_DOUT[0]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  10.62 0 10.88 0.26 ;
        END
    END A_DOUT[0]
    PIN A_ADDR[0]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 8.9011 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 45.2233 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  388.44 0 388.7 0.26 ;
        END
    END A_ADDR[0]
    PIN A_BIST_ADDR[0]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 9.6967 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 49.1845 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  393.03 0 393.29 0.26 ;
        END
    END A_BIST_ADDR[0]
    PIN A_ADDR[1]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 7.774 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 39.657 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  387.93 0 388.19 0.26 ;
        END
    END A_ADDR[1]
    PIN A_BIST_ADDR[1]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 8.5696 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 43.6181 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  392.52 0 392.78 0.26 ;
        END
    END A_BIST_ADDR[1]
    PIN A_ADDR[2]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 10.6327 LAYER Metal2 ;
        ANTENNAPARTIALMETALAREA 1.5246 LAYER Metal3 ;
        ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
        ANTENNAMAXAREACAR 9.41598 LAYER Metal3 ;
        PORT
            LAYER Metal2 ;
              RECT  396.09 0 396.35 0.26 ;
        END
    END A_ADDR[2]
    PIN A_BIST_ADDR[2]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 10.6327 LAYER Metal2 ;
        ANTENNAPARTIALMETALAREA 1.0962 LAYER Metal3 ;
        ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
        ANTENNAMAXAREACAR 7.81379 LAYER Metal3 ;
        PORT
            LAYER Metal2 ;
              RECT  396.6 0 396.86 0.26 ;
        END
    END A_BIST_ADDR[2]
    PIN A_ADDR[3]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 10.6327 LAYER Metal2 ;
        ANTENNAPARTIALMETALAREA 3.8367 LAYER Metal3 ;
        ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
        ANTENNAMAXAREACAR 20.9276 LAYER Metal3 ;
        PORT
            LAYER Metal2 ;
              RECT  395.07 0 395.33 0.26 ;
        END
    END A_ADDR[3]
    PIN A_BIST_ADDR[3]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 10.6327 LAYER Metal2 ;
        ANTENNAPARTIALMETALAREA 3.5175 LAYER Metal3 ;
        ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
        ANTENNAMAXAREACAR 19.8691 LAYER Metal3 ;
        PORT
            LAYER Metal2 ;
              RECT  395.58 0 395.84 0.26 ;
        END
    END A_BIST_ADDR[3]
    PIN A_ADDR[4]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 12.1979 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 61.6375 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  398.64 0 398.9 0.26 ;
        END
    END A_ADDR[4]
    PIN A_BIST_ADDR[4]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 11.9327 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 60.3172 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  398.13 0 398.39 0.26 ;
        END
    END A_BIST_ADDR[4]
    PIN A_ADDR[5]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 13.9269 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 70.246 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  397.62 0 397.88 0.26 ;
        END
    END A_ADDR[5]
    PIN A_BIST_ADDR[5]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 13.6617 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 68.9256 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  397.11 0 397.37 0.26 ;
        END
    END A_BIST_ADDR[5]
    PIN A_ADDR[6]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 10.9525 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 55.4369 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  376.2 0 376.46 0.26 ;
        END
    END A_ADDR[6]
    PIN A_BIST_ADDR[6]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 10.6771 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 54.0657 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  376.71 0 376.97 0.26 ;
        END
    END A_BIST_ADDR[6]
    PIN A_ADDR[7]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 12.4163 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 62.7249 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  377.22 0 377.48 0.26 ;
        END
    END A_ADDR[7]
    PIN A_BIST_ADDR[7]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 12.1511 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 61.4045 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  377.73 0 377.99 0.26 ;
        END
    END A_BIST_ADDR[7]
    PIN A_CLK
        DIRECTION INPUT ; 
        USE CLOCK ; 
        ANTENNAPARTIALMETALAREA 4.0547 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 21.0939 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  386.4 0 386.66 0.26 ;
        END
    END A_CLK
    PIN A_REN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.99505 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 20.7969 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  389.97 0 390.23 0.26 ;
        END
    END A_REN
    PIN A_WEN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 15.2686 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  389.46 0 389.72 0.26 ;
        END
    END A_WEN
    PIN A_MEN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.0247 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 15.9656 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  386.91 0 387.17 0.26 ;
        END
    END A_MEN
    PIN A_DLY
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 6.058 LAYER Metal2 ;
        ANTENNAGATEAREA 0.3367 LAYER Metal2 ;
        ANTENNAMAXAREACAR 18.5328 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  408.33 0 408.59 0.26 ;
        END
    END A_DLY
    PIN A_BIST_EN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.9871 LAYER Metal2 ;
        ANTENNAPARTIALMETALAREA 382.413 LAYER Metal3 ;
        ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
        ANTENNAGATEAREA 1.43 LAYER Metal2 ;
        ANTENNAGATEAREA 50.05 LAYER Metal3 ;
        ANTENNAMAXAREACAR 3.21364 LAYER Metal2 ;
        ANTENNAMAXAREACAR 17.9133 LAYER Metal3 ;
        ANTENNAMAXCUTCAR 0.151469 LAYER Via2 ;
        PORT
            LAYER Metal2 ;
              RECT  388.95 0 389.21 0.26 ;
        END
    END A_BIST_EN
    PIN A_BIST_CLK
        DIRECTION INPUT ; 
        USE CLOCK ; 
        ANTENNAPARTIALMETALAREA 4.1639 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 21.9534 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  384.87 0 385.13 0.26 ;
        END
    END A_BIST_CLK
    PIN A_BIST_REN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 4.1119 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 21.6945 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  391.5 0 391.76 0.26 ;
        END
    END A_BIST_REN
    PIN A_BIST_WEN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 2.9051 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 15.6861 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  390.99 0 391.25 0.26 ;
        END
    END A_BIST_WEN
    PIN A_BIST_MEN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 2.8977 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 15.6492 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  385.38 0 385.64 0.26 ;
        END
    END A_BIST_MEN
    OBS
      LAYER Metal1 ;
        RECT  0 0 784.48 118.78 ;
      LAYER Metal2 ;
        RECT  0.105 45.465 0.305 118.755 ;
        RECT  1.1 118.025 1.3 118.755 ;
        RECT  3.29 0.52 3.55 5.16 ;
        RECT  2.77 4.9 3.55 5.16 ;
        RECT  2.77 4.9 3.03 6.64 ;
        RECT  1.92 118.025 2.12 118.755 ;
        RECT  2.415 118.025 2.615 118.755 ;
        RECT  2.915 118.025 3.115 118.755 ;
        RECT  3.415 118.025 3.615 118.755 ;
        RECT  3.91 118.025 4.11 118.755 ;
        RECT  4.655 0.17 5.425 0.94 ;
        RECT  4.655 0.17 4.915 12.9 ;
        RECT  5.165 0.17 5.425 12.9 ;
        RECT  4.145 0.52 4.405 5.815 ;
        RECT  4.73 118.025 4.93 118.755 ;
        RECT  5.675 0.17 6.445 0.43 ;
        RECT  5.675 0.17 5.935 11.5 ;
        RECT  6.185 0.17 6.445 11.5 ;
        RECT  5.225 118.025 5.425 118.755 ;
        RECT  5.725 118.025 5.925 118.755 ;
        RECT  6.225 118.025 6.425 118.755 ;
        RECT  7.715 0.17 8.485 0.43 ;
        RECT  7.715 0.17 7.975 10.48 ;
        RECT  8.225 0.17 8.485 10.99 ;
        RECT  6.72 118.025 6.92 118.755 ;
        RECT  7.54 118.025 7.74 118.755 ;
        RECT  8.735 0.17 9.505 0.94 ;
        RECT  8.735 0.17 8.995 8.7 ;
        RECT  9.245 0.17 9.505 12.9 ;
        RECT  8.035 118.025 8.235 118.755 ;
        RECT  8.535 118.025 8.735 118.755 ;
        RECT  9.035 118.025 9.235 118.755 ;
        RECT  9.53 118.025 9.73 118.755 ;
        RECT  9.755 0.52 10.015 2.485 ;
        RECT  10.35 118.025 10.55 118.755 ;
        RECT  10.62 0.52 10.88 14.11 ;
        RECT  10.845 118.025 11.045 118.755 ;
        RECT  11.13 0.52 11.39 2.335 ;
        RECT  11.345 118.025 11.545 118.755 ;
        RECT  11.845 118.025 12.045 118.755 ;
        RECT  12.34 118.025 12.54 118.755 ;
        RECT  14.53 0.52 14.79 5.16 ;
        RECT  14.01 4.9 14.79 5.16 ;
        RECT  14.01 4.9 14.27 6.64 ;
        RECT  13.16 118.025 13.36 118.755 ;
        RECT  13.655 118.025 13.855 118.755 ;
        RECT  14.155 118.025 14.355 118.755 ;
        RECT  14.655 118.025 14.855 118.755 ;
        RECT  15.15 118.025 15.35 118.755 ;
        RECT  15.895 0.17 16.665 0.94 ;
        RECT  15.895 0.17 16.155 12.9 ;
        RECT  16.405 0.17 16.665 12.9 ;
        RECT  15.385 0.52 15.645 5.815 ;
        RECT  15.97 118.025 16.17 118.755 ;
        RECT  16.915 0.17 17.685 0.43 ;
        RECT  16.915 0.17 17.175 11.5 ;
        RECT  17.425 0.17 17.685 11.5 ;
        RECT  16.465 118.025 16.665 118.755 ;
        RECT  16.965 118.025 17.165 118.755 ;
        RECT  17.465 118.025 17.665 118.755 ;
        RECT  18.955 0.17 19.725 0.43 ;
        RECT  18.955 0.17 19.215 10.48 ;
        RECT  19.465 0.17 19.725 10.99 ;
        RECT  17.96 118.025 18.16 118.755 ;
        RECT  18.78 118.025 18.98 118.755 ;
        RECT  19.975 0.17 20.745 0.94 ;
        RECT  19.975 0.17 20.235 8.7 ;
        RECT  20.485 0.17 20.745 12.9 ;
        RECT  19.275 118.025 19.475 118.755 ;
        RECT  19.775 118.025 19.975 118.755 ;
        RECT  20.275 118.025 20.475 118.755 ;
        RECT  20.77 118.025 20.97 118.755 ;
        RECT  20.995 0.52 21.255 2.485 ;
        RECT  21.59 118.025 21.79 118.755 ;
        RECT  21.86 0.52 22.12 14.11 ;
        RECT  22.085 118.025 22.285 118.755 ;
        RECT  22.37 0.52 22.63 2.335 ;
        RECT  22.585 118.025 22.785 118.755 ;
        RECT  23.085 118.025 23.285 118.755 ;
        RECT  23.58 118.025 23.78 118.755 ;
        RECT  25.77 0.52 26.03 5.16 ;
        RECT  25.25 4.9 26.03 5.16 ;
        RECT  25.25 4.9 25.51 6.64 ;
        RECT  24.4 118.025 24.6 118.755 ;
        RECT  24.895 118.025 25.095 118.755 ;
        RECT  25.395 118.025 25.595 118.755 ;
        RECT  25.895 118.025 26.095 118.755 ;
        RECT  26.39 118.025 26.59 118.755 ;
        RECT  27.135 0.17 27.905 0.94 ;
        RECT  27.135 0.17 27.395 12.9 ;
        RECT  27.645 0.17 27.905 12.9 ;
        RECT  26.625 0.52 26.885 5.815 ;
        RECT  27.21 118.025 27.41 118.755 ;
        RECT  28.155 0.17 28.925 0.43 ;
        RECT  28.155 0.17 28.415 11.5 ;
        RECT  28.665 0.17 28.925 11.5 ;
        RECT  27.705 118.025 27.905 118.755 ;
        RECT  28.205 118.025 28.405 118.755 ;
        RECT  28.705 118.025 28.905 118.755 ;
        RECT  30.195 0.17 30.965 0.43 ;
        RECT  30.195 0.17 30.455 10.48 ;
        RECT  30.705 0.17 30.965 10.99 ;
        RECT  29.2 118.025 29.4 118.755 ;
        RECT  30.02 118.025 30.22 118.755 ;
        RECT  31.215 0.17 31.985 0.94 ;
        RECT  31.215 0.17 31.475 8.7 ;
        RECT  31.725 0.17 31.985 12.9 ;
        RECT  30.515 118.025 30.715 118.755 ;
        RECT  31.015 118.025 31.215 118.755 ;
        RECT  31.515 118.025 31.715 118.755 ;
        RECT  32.01 118.025 32.21 118.755 ;
        RECT  32.235 0.52 32.495 2.485 ;
        RECT  32.83 118.025 33.03 118.755 ;
        RECT  33.1 0.52 33.36 14.11 ;
        RECT  33.325 118.025 33.525 118.755 ;
        RECT  33.61 0.52 33.87 2.335 ;
        RECT  33.825 118.025 34.025 118.755 ;
        RECT  34.325 118.025 34.525 118.755 ;
        RECT  34.82 118.025 35.02 118.755 ;
        RECT  37.01 0.52 37.27 5.16 ;
        RECT  36.49 4.9 37.27 5.16 ;
        RECT  36.49 4.9 36.75 6.64 ;
        RECT  35.64 118.025 35.84 118.755 ;
        RECT  36.135 118.025 36.335 118.755 ;
        RECT  36.635 118.025 36.835 118.755 ;
        RECT  37.135 118.025 37.335 118.755 ;
        RECT  37.63 118.025 37.83 118.755 ;
        RECT  38.375 0.17 39.145 0.94 ;
        RECT  38.375 0.17 38.635 12.9 ;
        RECT  38.885 0.17 39.145 12.9 ;
        RECT  37.865 0.52 38.125 5.815 ;
        RECT  38.45 118.025 38.65 118.755 ;
        RECT  39.395 0.17 40.165 0.43 ;
        RECT  39.395 0.17 39.655 11.5 ;
        RECT  39.905 0.17 40.165 11.5 ;
        RECT  38.945 118.025 39.145 118.755 ;
        RECT  39.445 118.025 39.645 118.755 ;
        RECT  39.945 118.025 40.145 118.755 ;
        RECT  41.435 0.17 42.205 0.43 ;
        RECT  41.435 0.17 41.695 10.48 ;
        RECT  41.945 0.17 42.205 10.99 ;
        RECT  40.44 118.025 40.64 118.755 ;
        RECT  41.26 118.025 41.46 118.755 ;
        RECT  42.455 0.17 43.225 0.94 ;
        RECT  42.455 0.17 42.715 8.7 ;
        RECT  42.965 0.17 43.225 12.9 ;
        RECT  41.755 118.025 41.955 118.755 ;
        RECT  42.255 118.025 42.455 118.755 ;
        RECT  42.755 118.025 42.955 118.755 ;
        RECT  43.25 118.025 43.45 118.755 ;
        RECT  43.475 0.52 43.735 2.485 ;
        RECT  44.07 118.025 44.27 118.755 ;
        RECT  44.34 0.52 44.6 14.11 ;
        RECT  44.565 118.025 44.765 118.755 ;
        RECT  44.85 0.52 45.11 2.335 ;
        RECT  45.065 118.025 45.265 118.755 ;
        RECT  45.565 118.025 45.765 118.755 ;
        RECT  46.06 118.025 46.26 118.755 ;
        RECT  48.25 0.52 48.51 5.16 ;
        RECT  47.73 4.9 48.51 5.16 ;
        RECT  47.73 4.9 47.99 6.64 ;
        RECT  46.88 118.025 47.08 118.755 ;
        RECT  47.375 118.025 47.575 118.755 ;
        RECT  47.875 118.025 48.075 118.755 ;
        RECT  48.375 118.025 48.575 118.755 ;
        RECT  48.87 118.025 49.07 118.755 ;
        RECT  49.615 0.17 50.385 0.94 ;
        RECT  49.615 0.17 49.875 12.9 ;
        RECT  50.125 0.17 50.385 12.9 ;
        RECT  49.105 0.52 49.365 5.815 ;
        RECT  49.69 118.025 49.89 118.755 ;
        RECT  50.635 0.17 51.405 0.43 ;
        RECT  50.635 0.17 50.895 11.5 ;
        RECT  51.145 0.17 51.405 11.5 ;
        RECT  50.185 118.025 50.385 118.755 ;
        RECT  50.685 118.025 50.885 118.755 ;
        RECT  51.185 118.025 51.385 118.755 ;
        RECT  52.675 0.17 53.445 0.43 ;
        RECT  52.675 0.17 52.935 10.48 ;
        RECT  53.185 0.17 53.445 10.99 ;
        RECT  51.68 118.025 51.88 118.755 ;
        RECT  52.5 118.025 52.7 118.755 ;
        RECT  53.695 0.17 54.465 0.94 ;
        RECT  53.695 0.17 53.955 8.7 ;
        RECT  54.205 0.17 54.465 12.9 ;
        RECT  52.995 118.025 53.195 118.755 ;
        RECT  53.495 118.025 53.695 118.755 ;
        RECT  53.995 118.025 54.195 118.755 ;
        RECT  54.49 118.025 54.69 118.755 ;
        RECT  54.715 0.52 54.975 2.485 ;
        RECT  55.31 118.025 55.51 118.755 ;
        RECT  55.58 0.52 55.84 14.11 ;
        RECT  55.805 118.025 56.005 118.755 ;
        RECT  56.09 0.52 56.35 2.335 ;
        RECT  56.305 118.025 56.505 118.755 ;
        RECT  56.805 118.025 57.005 118.755 ;
        RECT  57.3 118.025 57.5 118.755 ;
        RECT  59.49 0.52 59.75 5.16 ;
        RECT  58.97 4.9 59.75 5.16 ;
        RECT  58.97 4.9 59.23 6.64 ;
        RECT  58.12 118.025 58.32 118.755 ;
        RECT  58.615 118.025 58.815 118.755 ;
        RECT  59.115 118.025 59.315 118.755 ;
        RECT  59.615 118.025 59.815 118.755 ;
        RECT  60.11 118.025 60.31 118.755 ;
        RECT  60.855 0.17 61.625 0.94 ;
        RECT  60.855 0.17 61.115 12.9 ;
        RECT  61.365 0.17 61.625 12.9 ;
        RECT  60.345 0.52 60.605 5.815 ;
        RECT  60.93 118.025 61.13 118.755 ;
        RECT  61.875 0.17 62.645 0.43 ;
        RECT  61.875 0.17 62.135 11.5 ;
        RECT  62.385 0.17 62.645 11.5 ;
        RECT  61.425 118.025 61.625 118.755 ;
        RECT  61.925 118.025 62.125 118.755 ;
        RECT  62.425 118.025 62.625 118.755 ;
        RECT  63.915 0.17 64.685 0.43 ;
        RECT  63.915 0.17 64.175 10.48 ;
        RECT  64.425 0.17 64.685 10.99 ;
        RECT  62.92 118.025 63.12 118.755 ;
        RECT  63.74 118.025 63.94 118.755 ;
        RECT  64.935 0.17 65.705 0.94 ;
        RECT  64.935 0.17 65.195 8.7 ;
        RECT  65.445 0.17 65.705 12.9 ;
        RECT  64.235 118.025 64.435 118.755 ;
        RECT  64.735 118.025 64.935 118.755 ;
        RECT  65.235 118.025 65.435 118.755 ;
        RECT  65.73 118.025 65.93 118.755 ;
        RECT  65.955 0.52 66.215 2.485 ;
        RECT  66.55 118.025 66.75 118.755 ;
        RECT  66.82 0.52 67.08 14.11 ;
        RECT  67.045 118.025 67.245 118.755 ;
        RECT  67.33 0.52 67.59 2.335 ;
        RECT  67.545 118.025 67.745 118.755 ;
        RECT  68.045 118.025 68.245 118.755 ;
        RECT  68.54 118.025 68.74 118.755 ;
        RECT  70.73 0.52 70.99 5.16 ;
        RECT  70.21 4.9 70.99 5.16 ;
        RECT  70.21 4.9 70.47 6.64 ;
        RECT  69.36 118.025 69.56 118.755 ;
        RECT  69.855 118.025 70.055 118.755 ;
        RECT  70.355 118.025 70.555 118.755 ;
        RECT  70.855 118.025 71.055 118.755 ;
        RECT  71.35 118.025 71.55 118.755 ;
        RECT  72.095 0.17 72.865 0.94 ;
        RECT  72.095 0.17 72.355 12.9 ;
        RECT  72.605 0.17 72.865 12.9 ;
        RECT  71.585 0.52 71.845 5.815 ;
        RECT  72.17 118.025 72.37 118.755 ;
        RECT  73.115 0.17 73.885 0.43 ;
        RECT  73.115 0.17 73.375 11.5 ;
        RECT  73.625 0.17 73.885 11.5 ;
        RECT  72.665 118.025 72.865 118.755 ;
        RECT  73.165 118.025 73.365 118.755 ;
        RECT  73.665 118.025 73.865 118.755 ;
        RECT  75.155 0.17 75.925 0.43 ;
        RECT  75.155 0.17 75.415 10.48 ;
        RECT  75.665 0.17 75.925 10.99 ;
        RECT  74.16 118.025 74.36 118.755 ;
        RECT  74.98 118.025 75.18 118.755 ;
        RECT  76.175 0.17 76.945 0.94 ;
        RECT  76.175 0.17 76.435 8.7 ;
        RECT  76.685 0.17 76.945 12.9 ;
        RECT  75.475 118.025 75.675 118.755 ;
        RECT  75.975 118.025 76.175 118.755 ;
        RECT  76.475 118.025 76.675 118.755 ;
        RECT  76.97 118.025 77.17 118.755 ;
        RECT  77.195 0.52 77.455 2.485 ;
        RECT  77.79 118.025 77.99 118.755 ;
        RECT  78.06 0.52 78.32 14.11 ;
        RECT  78.285 118.025 78.485 118.755 ;
        RECT  78.57 0.52 78.83 2.335 ;
        RECT  78.785 118.025 78.985 118.755 ;
        RECT  79.285 118.025 79.485 118.755 ;
        RECT  79.78 118.025 79.98 118.755 ;
        RECT  81.97 0.52 82.23 5.16 ;
        RECT  81.45 4.9 82.23 5.16 ;
        RECT  81.45 4.9 81.71 6.64 ;
        RECT  80.6 118.025 80.8 118.755 ;
        RECT  81.095 118.025 81.295 118.755 ;
        RECT  81.595 118.025 81.795 118.755 ;
        RECT  82.095 118.025 82.295 118.755 ;
        RECT  82.59 118.025 82.79 118.755 ;
        RECT  83.335 0.17 84.105 0.94 ;
        RECT  83.335 0.17 83.595 12.9 ;
        RECT  83.845 0.17 84.105 12.9 ;
        RECT  82.825 0.52 83.085 5.815 ;
        RECT  83.41 118.025 83.61 118.755 ;
        RECT  84.355 0.17 85.125 0.43 ;
        RECT  84.355 0.17 84.615 11.5 ;
        RECT  84.865 0.17 85.125 11.5 ;
        RECT  83.905 118.025 84.105 118.755 ;
        RECT  84.405 118.025 84.605 118.755 ;
        RECT  84.905 118.025 85.105 118.755 ;
        RECT  86.395 0.17 87.165 0.43 ;
        RECT  86.395 0.17 86.655 10.48 ;
        RECT  86.905 0.17 87.165 10.99 ;
        RECT  85.4 118.025 85.6 118.755 ;
        RECT  86.22 118.025 86.42 118.755 ;
        RECT  87.415 0.17 88.185 0.94 ;
        RECT  87.415 0.17 87.675 8.7 ;
        RECT  87.925 0.17 88.185 12.9 ;
        RECT  86.715 118.025 86.915 118.755 ;
        RECT  87.215 118.025 87.415 118.755 ;
        RECT  87.715 118.025 87.915 118.755 ;
        RECT  88.21 118.025 88.41 118.755 ;
        RECT  88.435 0.52 88.695 2.485 ;
        RECT  89.03 118.025 89.23 118.755 ;
        RECT  89.3 0.52 89.56 14.11 ;
        RECT  89.525 118.025 89.725 118.755 ;
        RECT  89.81 0.52 90.07 2.335 ;
        RECT  90.025 118.025 90.225 118.755 ;
        RECT  90.525 118.025 90.725 118.755 ;
        RECT  91.02 118.025 91.22 118.755 ;
        RECT  93.21 0.52 93.47 5.16 ;
        RECT  92.69 4.9 93.47 5.16 ;
        RECT  92.69 4.9 92.95 6.64 ;
        RECT  91.84 118.025 92.04 118.755 ;
        RECT  92.335 118.025 92.535 118.755 ;
        RECT  92.835 118.025 93.035 118.755 ;
        RECT  93.335 118.025 93.535 118.755 ;
        RECT  93.83 118.025 94.03 118.755 ;
        RECT  94.575 0.17 95.345 0.94 ;
        RECT  94.575 0.17 94.835 12.9 ;
        RECT  95.085 0.17 95.345 12.9 ;
        RECT  94.065 0.52 94.325 5.815 ;
        RECT  94.65 118.025 94.85 118.755 ;
        RECT  95.595 0.17 96.365 0.43 ;
        RECT  95.595 0.17 95.855 11.5 ;
        RECT  96.105 0.17 96.365 11.5 ;
        RECT  95.145 118.025 95.345 118.755 ;
        RECT  95.645 118.025 95.845 118.755 ;
        RECT  96.145 118.025 96.345 118.755 ;
        RECT  97.635 0.17 98.405 0.43 ;
        RECT  97.635 0.17 97.895 10.48 ;
        RECT  98.145 0.17 98.405 10.99 ;
        RECT  96.64 118.025 96.84 118.755 ;
        RECT  97.46 118.025 97.66 118.755 ;
        RECT  98.655 0.17 99.425 0.94 ;
        RECT  98.655 0.17 98.915 8.7 ;
        RECT  99.165 0.17 99.425 12.9 ;
        RECT  97.955 118.025 98.155 118.755 ;
        RECT  98.455 118.025 98.655 118.755 ;
        RECT  98.955 118.025 99.155 118.755 ;
        RECT  99.45 118.025 99.65 118.755 ;
        RECT  99.675 0.52 99.935 2.485 ;
        RECT  100.27 118.025 100.47 118.755 ;
        RECT  100.54 0.52 100.8 14.11 ;
        RECT  100.765 118.025 100.965 118.755 ;
        RECT  101.05 0.52 101.31 2.335 ;
        RECT  101.265 118.025 101.465 118.755 ;
        RECT  101.765 118.025 101.965 118.755 ;
        RECT  102.26 118.025 102.46 118.755 ;
        RECT  104.45 0.52 104.71 5.16 ;
        RECT  103.93 4.9 104.71 5.16 ;
        RECT  103.93 4.9 104.19 6.64 ;
        RECT  103.08 118.025 103.28 118.755 ;
        RECT  103.575 118.025 103.775 118.755 ;
        RECT  104.075 118.025 104.275 118.755 ;
        RECT  104.575 118.025 104.775 118.755 ;
        RECT  105.07 118.025 105.27 118.755 ;
        RECT  105.815 0.17 106.585 0.94 ;
        RECT  105.815 0.17 106.075 12.9 ;
        RECT  106.325 0.17 106.585 12.9 ;
        RECT  105.305 0.52 105.565 5.815 ;
        RECT  105.89 118.025 106.09 118.755 ;
        RECT  106.835 0.17 107.605 0.43 ;
        RECT  106.835 0.17 107.095 11.5 ;
        RECT  107.345 0.17 107.605 11.5 ;
        RECT  106.385 118.025 106.585 118.755 ;
        RECT  106.885 118.025 107.085 118.755 ;
        RECT  107.385 118.025 107.585 118.755 ;
        RECT  108.875 0.17 109.645 0.43 ;
        RECT  108.875 0.17 109.135 10.48 ;
        RECT  109.385 0.17 109.645 10.99 ;
        RECT  107.88 118.025 108.08 118.755 ;
        RECT  108.7 118.025 108.9 118.755 ;
        RECT  109.895 0.17 110.665 0.94 ;
        RECT  109.895 0.17 110.155 8.7 ;
        RECT  110.405 0.17 110.665 12.9 ;
        RECT  109.195 118.025 109.395 118.755 ;
        RECT  109.695 118.025 109.895 118.755 ;
        RECT  110.195 118.025 110.395 118.755 ;
        RECT  110.69 118.025 110.89 118.755 ;
        RECT  110.915 0.52 111.175 2.485 ;
        RECT  111.51 118.025 111.71 118.755 ;
        RECT  111.78 0.52 112.04 14.11 ;
        RECT  112.005 118.025 112.205 118.755 ;
        RECT  112.29 0.52 112.55 2.335 ;
        RECT  112.505 118.025 112.705 118.755 ;
        RECT  113.005 118.025 113.205 118.755 ;
        RECT  113.5 118.025 113.7 118.755 ;
        RECT  115.69 0.52 115.95 5.16 ;
        RECT  115.17 4.9 115.95 5.16 ;
        RECT  115.17 4.9 115.43 6.64 ;
        RECT  114.32 118.025 114.52 118.755 ;
        RECT  114.815 118.025 115.015 118.755 ;
        RECT  115.315 118.025 115.515 118.755 ;
        RECT  115.815 118.025 116.015 118.755 ;
        RECT  116.31 118.025 116.51 118.755 ;
        RECT  117.055 0.17 117.825 0.94 ;
        RECT  117.055 0.17 117.315 12.9 ;
        RECT  117.565 0.17 117.825 12.9 ;
        RECT  116.545 0.52 116.805 5.815 ;
        RECT  117.13 118.025 117.33 118.755 ;
        RECT  118.075 0.17 118.845 0.43 ;
        RECT  118.075 0.17 118.335 11.5 ;
        RECT  118.585 0.17 118.845 11.5 ;
        RECT  117.625 118.025 117.825 118.755 ;
        RECT  118.125 118.025 118.325 118.755 ;
        RECT  118.625 118.025 118.825 118.755 ;
        RECT  120.115 0.17 120.885 0.43 ;
        RECT  120.115 0.17 120.375 10.48 ;
        RECT  120.625 0.17 120.885 10.99 ;
        RECT  119.12 118.025 119.32 118.755 ;
        RECT  119.94 118.025 120.14 118.755 ;
        RECT  121.135 0.17 121.905 0.94 ;
        RECT  121.135 0.17 121.395 8.7 ;
        RECT  121.645 0.17 121.905 12.9 ;
        RECT  120.435 118.025 120.635 118.755 ;
        RECT  120.935 118.025 121.135 118.755 ;
        RECT  121.435 118.025 121.635 118.755 ;
        RECT  121.93 118.025 122.13 118.755 ;
        RECT  122.155 0.52 122.415 2.485 ;
        RECT  122.75 118.025 122.95 118.755 ;
        RECT  123.02 0.52 123.28 14.11 ;
        RECT  123.245 118.025 123.445 118.755 ;
        RECT  123.53 0.52 123.79 2.335 ;
        RECT  123.745 118.025 123.945 118.755 ;
        RECT  124.245 118.025 124.445 118.755 ;
        RECT  124.74 118.025 124.94 118.755 ;
        RECT  126.93 0.52 127.19 5.16 ;
        RECT  126.41 4.9 127.19 5.16 ;
        RECT  126.41 4.9 126.67 6.64 ;
        RECT  125.56 118.025 125.76 118.755 ;
        RECT  126.055 118.025 126.255 118.755 ;
        RECT  126.555 118.025 126.755 118.755 ;
        RECT  127.055 118.025 127.255 118.755 ;
        RECT  127.55 118.025 127.75 118.755 ;
        RECT  128.295 0.17 129.065 0.94 ;
        RECT  128.295 0.17 128.555 12.9 ;
        RECT  128.805 0.17 129.065 12.9 ;
        RECT  127.785 0.52 128.045 5.815 ;
        RECT  128.37 118.025 128.57 118.755 ;
        RECT  129.315 0.17 130.085 0.43 ;
        RECT  129.315 0.17 129.575 11.5 ;
        RECT  129.825 0.17 130.085 11.5 ;
        RECT  128.865 118.025 129.065 118.755 ;
        RECT  129.365 118.025 129.565 118.755 ;
        RECT  129.865 118.025 130.065 118.755 ;
        RECT  131.355 0.17 132.125 0.43 ;
        RECT  131.355 0.17 131.615 10.48 ;
        RECT  131.865 0.17 132.125 10.99 ;
        RECT  130.36 118.025 130.56 118.755 ;
        RECT  131.18 118.025 131.38 118.755 ;
        RECT  132.375 0.17 133.145 0.94 ;
        RECT  132.375 0.17 132.635 8.7 ;
        RECT  132.885 0.17 133.145 12.9 ;
        RECT  131.675 118.025 131.875 118.755 ;
        RECT  132.175 118.025 132.375 118.755 ;
        RECT  132.675 118.025 132.875 118.755 ;
        RECT  133.17 118.025 133.37 118.755 ;
        RECT  133.395 0.52 133.655 2.485 ;
        RECT  133.99 118.025 134.19 118.755 ;
        RECT  134.26 0.52 134.52 14.11 ;
        RECT  134.485 118.025 134.685 118.755 ;
        RECT  134.77 0.52 135.03 2.335 ;
        RECT  134.985 118.025 135.185 118.755 ;
        RECT  135.485 118.025 135.685 118.755 ;
        RECT  135.98 118.025 136.18 118.755 ;
        RECT  138.17 0.52 138.43 5.16 ;
        RECT  137.65 4.9 138.43 5.16 ;
        RECT  137.65 4.9 137.91 6.64 ;
        RECT  136.8 118.025 137 118.755 ;
        RECT  137.295 118.025 137.495 118.755 ;
        RECT  137.795 118.025 137.995 118.755 ;
        RECT  138.295 118.025 138.495 118.755 ;
        RECT  138.79 118.025 138.99 118.755 ;
        RECT  139.535 0.17 140.305 0.94 ;
        RECT  139.535 0.17 139.795 12.9 ;
        RECT  140.045 0.17 140.305 12.9 ;
        RECT  139.025 0.52 139.285 5.815 ;
        RECT  139.61 118.025 139.81 118.755 ;
        RECT  140.555 0.17 141.325 0.43 ;
        RECT  140.555 0.17 140.815 11.5 ;
        RECT  141.065 0.17 141.325 11.5 ;
        RECT  140.105 118.025 140.305 118.755 ;
        RECT  140.605 118.025 140.805 118.755 ;
        RECT  141.105 118.025 141.305 118.755 ;
        RECT  142.595 0.17 143.365 0.43 ;
        RECT  142.595 0.17 142.855 10.48 ;
        RECT  143.105 0.17 143.365 10.99 ;
        RECT  141.6 118.025 141.8 118.755 ;
        RECT  142.42 118.025 142.62 118.755 ;
        RECT  143.615 0.17 144.385 0.94 ;
        RECT  143.615 0.17 143.875 8.7 ;
        RECT  144.125 0.17 144.385 12.9 ;
        RECT  142.915 118.025 143.115 118.755 ;
        RECT  143.415 118.025 143.615 118.755 ;
        RECT  143.915 118.025 144.115 118.755 ;
        RECT  144.41 118.025 144.61 118.755 ;
        RECT  144.635 0.52 144.895 2.485 ;
        RECT  145.23 118.025 145.43 118.755 ;
        RECT  145.5 0.52 145.76 14.11 ;
        RECT  145.725 118.025 145.925 118.755 ;
        RECT  146.01 0.52 146.27 2.335 ;
        RECT  146.225 118.025 146.425 118.755 ;
        RECT  146.725 118.025 146.925 118.755 ;
        RECT  147.22 118.025 147.42 118.755 ;
        RECT  149.41 0.52 149.67 5.16 ;
        RECT  148.89 4.9 149.67 5.16 ;
        RECT  148.89 4.9 149.15 6.64 ;
        RECT  148.04 118.025 148.24 118.755 ;
        RECT  148.535 118.025 148.735 118.755 ;
        RECT  149.035 118.025 149.235 118.755 ;
        RECT  149.535 118.025 149.735 118.755 ;
        RECT  150.03 118.025 150.23 118.755 ;
        RECT  150.775 0.17 151.545 0.94 ;
        RECT  150.775 0.17 151.035 12.9 ;
        RECT  151.285 0.17 151.545 12.9 ;
        RECT  150.265 0.52 150.525 5.815 ;
        RECT  150.85 118.025 151.05 118.755 ;
        RECT  151.795 0.17 152.565 0.43 ;
        RECT  151.795 0.17 152.055 11.5 ;
        RECT  152.305 0.17 152.565 11.5 ;
        RECT  151.345 118.025 151.545 118.755 ;
        RECT  151.845 118.025 152.045 118.755 ;
        RECT  152.345 118.025 152.545 118.755 ;
        RECT  153.835 0.17 154.605 0.43 ;
        RECT  153.835 0.17 154.095 10.48 ;
        RECT  154.345 0.17 154.605 10.99 ;
        RECT  152.84 118.025 153.04 118.755 ;
        RECT  153.66 118.025 153.86 118.755 ;
        RECT  154.855 0.17 155.625 0.94 ;
        RECT  154.855 0.17 155.115 8.7 ;
        RECT  155.365 0.17 155.625 12.9 ;
        RECT  154.155 118.025 154.355 118.755 ;
        RECT  154.655 118.025 154.855 118.755 ;
        RECT  155.155 118.025 155.355 118.755 ;
        RECT  155.65 118.025 155.85 118.755 ;
        RECT  155.875 0.52 156.135 2.485 ;
        RECT  156.47 118.025 156.67 118.755 ;
        RECT  156.74 0.52 157 14.11 ;
        RECT  156.965 118.025 157.165 118.755 ;
        RECT  157.25 0.52 157.51 2.335 ;
        RECT  157.465 118.025 157.665 118.755 ;
        RECT  157.965 118.025 158.165 118.755 ;
        RECT  158.46 118.025 158.66 118.755 ;
        RECT  160.65 0.52 160.91 5.16 ;
        RECT  160.13 4.9 160.91 5.16 ;
        RECT  160.13 4.9 160.39 6.64 ;
        RECT  159.28 118.025 159.48 118.755 ;
        RECT  159.775 118.025 159.975 118.755 ;
        RECT  160.275 118.025 160.475 118.755 ;
        RECT  160.775 118.025 160.975 118.755 ;
        RECT  161.27 118.025 161.47 118.755 ;
        RECT  162.015 0.17 162.785 0.94 ;
        RECT  162.015 0.17 162.275 12.9 ;
        RECT  162.525 0.17 162.785 12.9 ;
        RECT  161.505 0.52 161.765 5.815 ;
        RECT  162.09 118.025 162.29 118.755 ;
        RECT  163.035 0.17 163.805 0.43 ;
        RECT  163.035 0.17 163.295 11.5 ;
        RECT  163.545 0.17 163.805 11.5 ;
        RECT  162.585 118.025 162.785 118.755 ;
        RECT  163.085 118.025 163.285 118.755 ;
        RECT  163.585 118.025 163.785 118.755 ;
        RECT  165.075 0.17 165.845 0.43 ;
        RECT  165.075 0.17 165.335 10.48 ;
        RECT  165.585 0.17 165.845 10.99 ;
        RECT  164.08 118.025 164.28 118.755 ;
        RECT  164.9 118.025 165.1 118.755 ;
        RECT  166.095 0.17 166.865 0.94 ;
        RECT  166.095 0.17 166.355 8.7 ;
        RECT  166.605 0.17 166.865 12.9 ;
        RECT  165.395 118.025 165.595 118.755 ;
        RECT  165.895 118.025 166.095 118.755 ;
        RECT  166.395 118.025 166.595 118.755 ;
        RECT  166.89 118.025 167.09 118.755 ;
        RECT  167.115 0.52 167.375 2.485 ;
        RECT  167.71 118.025 167.91 118.755 ;
        RECT  167.98 0.52 168.24 14.11 ;
        RECT  168.205 118.025 168.405 118.755 ;
        RECT  168.49 0.52 168.75 2.335 ;
        RECT  168.705 118.025 168.905 118.755 ;
        RECT  169.205 118.025 169.405 118.755 ;
        RECT  169.7 118.025 169.9 118.755 ;
        RECT  171.89 0.52 172.15 5.16 ;
        RECT  171.37 4.9 172.15 5.16 ;
        RECT  171.37 4.9 171.63 6.64 ;
        RECT  170.52 118.025 170.72 118.755 ;
        RECT  171.015 118.025 171.215 118.755 ;
        RECT  171.515 118.025 171.715 118.755 ;
        RECT  172.015 118.025 172.215 118.755 ;
        RECT  172.51 118.025 172.71 118.755 ;
        RECT  173.255 0.17 174.025 0.94 ;
        RECT  173.255 0.17 173.515 12.9 ;
        RECT  173.765 0.17 174.025 12.9 ;
        RECT  172.745 0.52 173.005 5.815 ;
        RECT  173.33 118.025 173.53 118.755 ;
        RECT  174.275 0.17 175.045 0.43 ;
        RECT  174.275 0.17 174.535 11.5 ;
        RECT  174.785 0.17 175.045 11.5 ;
        RECT  173.825 118.025 174.025 118.755 ;
        RECT  174.325 118.025 174.525 118.755 ;
        RECT  174.825 118.025 175.025 118.755 ;
        RECT  176.315 0.17 177.085 0.43 ;
        RECT  176.315 0.17 176.575 10.48 ;
        RECT  176.825 0.17 177.085 10.99 ;
        RECT  175.32 118.025 175.52 118.755 ;
        RECT  176.14 118.025 176.34 118.755 ;
        RECT  177.335 0.17 178.105 0.94 ;
        RECT  177.335 0.17 177.595 8.7 ;
        RECT  177.845 0.17 178.105 12.9 ;
        RECT  176.635 118.025 176.835 118.755 ;
        RECT  177.135 118.025 177.335 118.755 ;
        RECT  177.635 118.025 177.835 118.755 ;
        RECT  178.13 118.025 178.33 118.755 ;
        RECT  178.355 0.52 178.615 2.485 ;
        RECT  178.95 118.025 179.15 118.755 ;
        RECT  179.22 0.52 179.48 14.11 ;
        RECT  179.445 118.025 179.645 118.755 ;
        RECT  179.73 0.52 179.99 2.335 ;
        RECT  179.945 118.025 180.145 118.755 ;
        RECT  180.445 118.025 180.645 118.755 ;
        RECT  180.94 118.025 181.14 118.755 ;
        RECT  183.13 0.52 183.39 5.16 ;
        RECT  182.61 4.9 183.39 5.16 ;
        RECT  182.61 4.9 182.87 6.64 ;
        RECT  181.76 118.025 181.96 118.755 ;
        RECT  182.255 118.025 182.455 118.755 ;
        RECT  182.755 118.025 182.955 118.755 ;
        RECT  183.255 118.025 183.455 118.755 ;
        RECT  183.75 118.025 183.95 118.755 ;
        RECT  184.495 0.17 185.265 0.94 ;
        RECT  184.495 0.17 184.755 12.9 ;
        RECT  185.005 0.17 185.265 12.9 ;
        RECT  183.985 0.52 184.245 5.815 ;
        RECT  184.57 118.025 184.77 118.755 ;
        RECT  185.515 0.17 186.285 0.43 ;
        RECT  185.515 0.17 185.775 11.5 ;
        RECT  186.025 0.17 186.285 11.5 ;
        RECT  185.065 118.025 185.265 118.755 ;
        RECT  185.565 118.025 185.765 118.755 ;
        RECT  186.065 118.025 186.265 118.755 ;
        RECT  187.555 0.17 188.325 0.43 ;
        RECT  187.555 0.17 187.815 10.48 ;
        RECT  188.065 0.17 188.325 10.99 ;
        RECT  186.56 118.025 186.76 118.755 ;
        RECT  187.38 118.025 187.58 118.755 ;
        RECT  188.575 0.17 189.345 0.94 ;
        RECT  188.575 0.17 188.835 8.7 ;
        RECT  189.085 0.17 189.345 12.9 ;
        RECT  187.875 118.025 188.075 118.755 ;
        RECT  188.375 118.025 188.575 118.755 ;
        RECT  188.875 118.025 189.075 118.755 ;
        RECT  189.37 118.025 189.57 118.755 ;
        RECT  189.595 0.52 189.855 2.485 ;
        RECT  190.19 118.025 190.39 118.755 ;
        RECT  190.46 0.52 190.72 14.11 ;
        RECT  190.685 118.025 190.885 118.755 ;
        RECT  190.97 0.52 191.23 2.335 ;
        RECT  191.185 118.025 191.385 118.755 ;
        RECT  191.685 118.025 191.885 118.755 ;
        RECT  192.18 118.025 192.38 118.755 ;
        RECT  194.37 0.52 194.63 5.16 ;
        RECT  193.85 4.9 194.63 5.16 ;
        RECT  193.85 4.9 194.11 6.64 ;
        RECT  193 118.025 193.2 118.755 ;
        RECT  193.495 118.025 193.695 118.755 ;
        RECT  193.995 118.025 194.195 118.755 ;
        RECT  194.495 118.025 194.695 118.755 ;
        RECT  194.99 118.025 195.19 118.755 ;
        RECT  195.735 0.17 196.505 0.94 ;
        RECT  195.735 0.17 195.995 12.9 ;
        RECT  196.245 0.17 196.505 12.9 ;
        RECT  195.225 0.52 195.485 5.815 ;
        RECT  195.81 118.025 196.01 118.755 ;
        RECT  196.755 0.17 197.525 0.43 ;
        RECT  196.755 0.17 197.015 11.5 ;
        RECT  197.265 0.17 197.525 11.5 ;
        RECT  196.305 118.025 196.505 118.755 ;
        RECT  196.805 118.025 197.005 118.755 ;
        RECT  197.305 118.025 197.505 118.755 ;
        RECT  198.795 0.17 199.565 0.43 ;
        RECT  198.795 0.17 199.055 10.48 ;
        RECT  199.305 0.17 199.565 10.99 ;
        RECT  197.8 118.025 198 118.755 ;
        RECT  198.62 118.025 198.82 118.755 ;
        RECT  199.815 0.17 200.585 0.94 ;
        RECT  199.815 0.17 200.075 8.7 ;
        RECT  200.325 0.17 200.585 12.9 ;
        RECT  199.115 118.025 199.315 118.755 ;
        RECT  199.615 118.025 199.815 118.755 ;
        RECT  200.115 118.025 200.315 118.755 ;
        RECT  200.61 118.025 200.81 118.755 ;
        RECT  200.835 0.52 201.095 2.485 ;
        RECT  201.43 118.025 201.63 118.755 ;
        RECT  201.7 0.52 201.96 14.11 ;
        RECT  201.925 118.025 202.125 118.755 ;
        RECT  202.21 0.52 202.47 2.335 ;
        RECT  202.425 118.025 202.625 118.755 ;
        RECT  202.925 118.025 203.125 118.755 ;
        RECT  203.42 118.025 203.62 118.755 ;
        RECT  205.61 0.52 205.87 5.16 ;
        RECT  205.09 4.9 205.87 5.16 ;
        RECT  205.09 4.9 205.35 6.64 ;
        RECT  204.24 118.025 204.44 118.755 ;
        RECT  204.735 118.025 204.935 118.755 ;
        RECT  205.235 118.025 205.435 118.755 ;
        RECT  205.735 118.025 205.935 118.755 ;
        RECT  206.23 118.025 206.43 118.755 ;
        RECT  206.975 0.17 207.745 0.94 ;
        RECT  206.975 0.17 207.235 12.9 ;
        RECT  207.485 0.17 207.745 12.9 ;
        RECT  206.465 0.52 206.725 5.815 ;
        RECT  207.05 118.025 207.25 118.755 ;
        RECT  207.995 0.17 208.765 0.43 ;
        RECT  207.995 0.17 208.255 11.5 ;
        RECT  208.505 0.17 208.765 11.5 ;
        RECT  207.545 118.025 207.745 118.755 ;
        RECT  208.045 118.025 208.245 118.755 ;
        RECT  208.545 118.025 208.745 118.755 ;
        RECT  210.035 0.17 210.805 0.43 ;
        RECT  210.035 0.17 210.295 10.48 ;
        RECT  210.545 0.17 210.805 10.99 ;
        RECT  209.04 118.025 209.24 118.755 ;
        RECT  209.86 118.025 210.06 118.755 ;
        RECT  211.055 0.17 211.825 0.94 ;
        RECT  211.055 0.17 211.315 8.7 ;
        RECT  211.565 0.17 211.825 12.9 ;
        RECT  210.355 118.025 210.555 118.755 ;
        RECT  210.855 118.025 211.055 118.755 ;
        RECT  211.355 118.025 211.555 118.755 ;
        RECT  211.85 118.025 212.05 118.755 ;
        RECT  212.075 0.52 212.335 2.485 ;
        RECT  212.67 118.025 212.87 118.755 ;
        RECT  212.94 0.52 213.2 14.11 ;
        RECT  213.165 118.025 213.365 118.755 ;
        RECT  213.45 0.52 213.71 2.335 ;
        RECT  213.665 118.025 213.865 118.755 ;
        RECT  214.165 118.025 214.365 118.755 ;
        RECT  214.66 118.025 214.86 118.755 ;
        RECT  216.85 0.52 217.11 5.16 ;
        RECT  216.33 4.9 217.11 5.16 ;
        RECT  216.33 4.9 216.59 6.64 ;
        RECT  215.48 118.025 215.68 118.755 ;
        RECT  215.975 118.025 216.175 118.755 ;
        RECT  216.475 118.025 216.675 118.755 ;
        RECT  216.975 118.025 217.175 118.755 ;
        RECT  217.47 118.025 217.67 118.755 ;
        RECT  218.215 0.17 218.985 0.94 ;
        RECT  218.215 0.17 218.475 12.9 ;
        RECT  218.725 0.17 218.985 12.9 ;
        RECT  217.705 0.52 217.965 5.815 ;
        RECT  218.29 118.025 218.49 118.755 ;
        RECT  219.235 0.17 220.005 0.43 ;
        RECT  219.235 0.17 219.495 11.5 ;
        RECT  219.745 0.17 220.005 11.5 ;
        RECT  218.785 118.025 218.985 118.755 ;
        RECT  219.285 118.025 219.485 118.755 ;
        RECT  219.785 118.025 219.985 118.755 ;
        RECT  221.275 0.17 222.045 0.43 ;
        RECT  221.275 0.17 221.535 10.48 ;
        RECT  221.785 0.17 222.045 10.99 ;
        RECT  220.28 118.025 220.48 118.755 ;
        RECT  221.1 118.025 221.3 118.755 ;
        RECT  222.295 0.17 223.065 0.94 ;
        RECT  222.295 0.17 222.555 8.7 ;
        RECT  222.805 0.17 223.065 12.9 ;
        RECT  221.595 118.025 221.795 118.755 ;
        RECT  222.095 118.025 222.295 118.755 ;
        RECT  222.595 118.025 222.795 118.755 ;
        RECT  223.09 118.025 223.29 118.755 ;
        RECT  223.315 0.52 223.575 2.485 ;
        RECT  223.91 118.025 224.11 118.755 ;
        RECT  224.18 0.52 224.44 14.11 ;
        RECT  224.405 118.025 224.605 118.755 ;
        RECT  224.69 0.52 224.95 2.335 ;
        RECT  224.905 118.025 225.105 118.755 ;
        RECT  225.405 118.025 225.605 118.755 ;
        RECT  225.9 118.025 226.1 118.755 ;
        RECT  228.09 0.52 228.35 5.16 ;
        RECT  227.57 4.9 228.35 5.16 ;
        RECT  227.57 4.9 227.83 6.64 ;
        RECT  226.72 118.025 226.92 118.755 ;
        RECT  227.215 118.025 227.415 118.755 ;
        RECT  227.715 118.025 227.915 118.755 ;
        RECT  228.215 118.025 228.415 118.755 ;
        RECT  228.71 118.025 228.91 118.755 ;
        RECT  229.455 0.17 230.225 0.94 ;
        RECT  229.455 0.17 229.715 12.9 ;
        RECT  229.965 0.17 230.225 12.9 ;
        RECT  228.945 0.52 229.205 5.815 ;
        RECT  229.53 118.025 229.73 118.755 ;
        RECT  230.475 0.17 231.245 0.43 ;
        RECT  230.475 0.17 230.735 11.5 ;
        RECT  230.985 0.17 231.245 11.5 ;
        RECT  230.025 118.025 230.225 118.755 ;
        RECT  230.525 118.025 230.725 118.755 ;
        RECT  231.025 118.025 231.225 118.755 ;
        RECT  232.515 0.17 233.285 0.43 ;
        RECT  232.515 0.17 232.775 10.48 ;
        RECT  233.025 0.17 233.285 10.99 ;
        RECT  231.52 118.025 231.72 118.755 ;
        RECT  232.34 118.025 232.54 118.755 ;
        RECT  233.535 0.17 234.305 0.94 ;
        RECT  233.535 0.17 233.795 8.7 ;
        RECT  234.045 0.17 234.305 12.9 ;
        RECT  232.835 118.025 233.035 118.755 ;
        RECT  233.335 118.025 233.535 118.755 ;
        RECT  233.835 118.025 234.035 118.755 ;
        RECT  234.33 118.025 234.53 118.755 ;
        RECT  234.555 0.52 234.815 2.485 ;
        RECT  235.15 118.025 235.35 118.755 ;
        RECT  235.42 0.52 235.68 14.11 ;
        RECT  235.645 118.025 235.845 118.755 ;
        RECT  235.93 0.52 236.19 2.335 ;
        RECT  236.145 118.025 236.345 118.755 ;
        RECT  236.645 118.025 236.845 118.755 ;
        RECT  237.14 118.025 237.34 118.755 ;
        RECT  239.33 0.52 239.59 5.16 ;
        RECT  238.81 4.9 239.59 5.16 ;
        RECT  238.81 4.9 239.07 6.64 ;
        RECT  237.96 118.025 238.16 118.755 ;
        RECT  238.455 118.025 238.655 118.755 ;
        RECT  238.955 118.025 239.155 118.755 ;
        RECT  239.455 118.025 239.655 118.755 ;
        RECT  239.95 118.025 240.15 118.755 ;
        RECT  240.695 0.17 241.465 0.94 ;
        RECT  240.695 0.17 240.955 12.9 ;
        RECT  241.205 0.17 241.465 12.9 ;
        RECT  240.185 0.52 240.445 5.815 ;
        RECT  240.77 118.025 240.97 118.755 ;
        RECT  241.715 0.17 242.485 0.43 ;
        RECT  241.715 0.17 241.975 11.5 ;
        RECT  242.225 0.17 242.485 11.5 ;
        RECT  241.265 118.025 241.465 118.755 ;
        RECT  241.765 118.025 241.965 118.755 ;
        RECT  242.265 118.025 242.465 118.755 ;
        RECT  243.755 0.17 244.525 0.43 ;
        RECT  243.755 0.17 244.015 10.48 ;
        RECT  244.265 0.17 244.525 10.99 ;
        RECT  242.76 118.025 242.96 118.755 ;
        RECT  243.58 118.025 243.78 118.755 ;
        RECT  244.775 0.17 245.545 0.94 ;
        RECT  244.775 0.17 245.035 8.7 ;
        RECT  245.285 0.17 245.545 12.9 ;
        RECT  244.075 118.025 244.275 118.755 ;
        RECT  244.575 118.025 244.775 118.755 ;
        RECT  245.075 118.025 245.275 118.755 ;
        RECT  245.57 118.025 245.77 118.755 ;
        RECT  245.795 0.52 246.055 2.485 ;
        RECT  246.39 118.025 246.59 118.755 ;
        RECT  246.66 0.52 246.92 14.11 ;
        RECT  246.885 118.025 247.085 118.755 ;
        RECT  247.17 0.52 247.43 2.335 ;
        RECT  247.385 118.025 247.585 118.755 ;
        RECT  247.885 118.025 248.085 118.755 ;
        RECT  248.38 118.025 248.58 118.755 ;
        RECT  250.57 0.52 250.83 5.16 ;
        RECT  250.05 4.9 250.83 5.16 ;
        RECT  250.05 4.9 250.31 6.64 ;
        RECT  249.2 118.025 249.4 118.755 ;
        RECT  249.695 118.025 249.895 118.755 ;
        RECT  250.195 118.025 250.395 118.755 ;
        RECT  250.695 118.025 250.895 118.755 ;
        RECT  251.19 118.025 251.39 118.755 ;
        RECT  251.935 0.17 252.705 0.94 ;
        RECT  251.935 0.17 252.195 12.9 ;
        RECT  252.445 0.17 252.705 12.9 ;
        RECT  251.425 0.52 251.685 5.815 ;
        RECT  252.01 118.025 252.21 118.755 ;
        RECT  252.955 0.17 253.725 0.43 ;
        RECT  252.955 0.17 253.215 11.5 ;
        RECT  253.465 0.17 253.725 11.5 ;
        RECT  252.505 118.025 252.705 118.755 ;
        RECT  253.005 118.025 253.205 118.755 ;
        RECT  253.505 118.025 253.705 118.755 ;
        RECT  254.995 0.17 255.765 0.43 ;
        RECT  254.995 0.17 255.255 10.48 ;
        RECT  255.505 0.17 255.765 10.99 ;
        RECT  254 118.025 254.2 118.755 ;
        RECT  254.82 118.025 255.02 118.755 ;
        RECT  256.015 0.17 256.785 0.94 ;
        RECT  256.015 0.17 256.275 8.7 ;
        RECT  256.525 0.17 256.785 12.9 ;
        RECT  255.315 118.025 255.515 118.755 ;
        RECT  255.815 118.025 256.015 118.755 ;
        RECT  256.315 118.025 256.515 118.755 ;
        RECT  256.81 118.025 257.01 118.755 ;
        RECT  257.035 0.52 257.295 2.485 ;
        RECT  257.63 118.025 257.83 118.755 ;
        RECT  257.9 0.52 258.16 14.11 ;
        RECT  258.125 118.025 258.325 118.755 ;
        RECT  258.41 0.52 258.67 2.335 ;
        RECT  258.625 118.025 258.825 118.755 ;
        RECT  259.125 118.025 259.325 118.755 ;
        RECT  259.62 118.025 259.82 118.755 ;
        RECT  261.81 0.52 262.07 5.16 ;
        RECT  261.29 4.9 262.07 5.16 ;
        RECT  261.29 4.9 261.55 6.64 ;
        RECT  260.44 118.025 260.64 118.755 ;
        RECT  260.935 118.025 261.135 118.755 ;
        RECT  261.435 118.025 261.635 118.755 ;
        RECT  261.935 118.025 262.135 118.755 ;
        RECT  262.43 118.025 262.63 118.755 ;
        RECT  263.175 0.17 263.945 0.94 ;
        RECT  263.175 0.17 263.435 12.9 ;
        RECT  263.685 0.17 263.945 12.9 ;
        RECT  262.665 0.52 262.925 5.815 ;
        RECT  263.25 118.025 263.45 118.755 ;
        RECT  264.195 0.17 264.965 0.43 ;
        RECT  264.195 0.17 264.455 11.5 ;
        RECT  264.705 0.17 264.965 11.5 ;
        RECT  263.745 118.025 263.945 118.755 ;
        RECT  264.245 118.025 264.445 118.755 ;
        RECT  264.745 118.025 264.945 118.755 ;
        RECT  266.235 0.17 267.005 0.43 ;
        RECT  266.235 0.17 266.495 10.48 ;
        RECT  266.745 0.17 267.005 10.99 ;
        RECT  265.24 118.025 265.44 118.755 ;
        RECT  266.06 118.025 266.26 118.755 ;
        RECT  267.255 0.17 268.025 0.94 ;
        RECT  267.255 0.17 267.515 8.7 ;
        RECT  267.765 0.17 268.025 12.9 ;
        RECT  266.555 118.025 266.755 118.755 ;
        RECT  267.055 118.025 267.255 118.755 ;
        RECT  267.555 118.025 267.755 118.755 ;
        RECT  268.05 118.025 268.25 118.755 ;
        RECT  268.275 0.52 268.535 2.485 ;
        RECT  268.87 118.025 269.07 118.755 ;
        RECT  269.14 0.52 269.4 14.11 ;
        RECT  269.365 118.025 269.565 118.755 ;
        RECT  269.65 0.52 269.91 2.335 ;
        RECT  269.865 118.025 270.065 118.755 ;
        RECT  270.365 118.025 270.565 118.755 ;
        RECT  270.86 118.025 271.06 118.755 ;
        RECT  273.05 0.52 273.31 5.16 ;
        RECT  272.53 4.9 273.31 5.16 ;
        RECT  272.53 4.9 272.79 6.64 ;
        RECT  271.68 118.025 271.88 118.755 ;
        RECT  272.175 118.025 272.375 118.755 ;
        RECT  272.675 118.025 272.875 118.755 ;
        RECT  273.175 118.025 273.375 118.755 ;
        RECT  273.67 118.025 273.87 118.755 ;
        RECT  274.415 0.17 275.185 0.94 ;
        RECT  274.415 0.17 274.675 12.9 ;
        RECT  274.925 0.17 275.185 12.9 ;
        RECT  273.905 0.52 274.165 5.815 ;
        RECT  274.49 118.025 274.69 118.755 ;
        RECT  275.435 0.17 276.205 0.43 ;
        RECT  275.435 0.17 275.695 11.5 ;
        RECT  275.945 0.17 276.205 11.5 ;
        RECT  274.985 118.025 275.185 118.755 ;
        RECT  275.485 118.025 275.685 118.755 ;
        RECT  275.985 118.025 276.185 118.755 ;
        RECT  277.475 0.17 278.245 0.43 ;
        RECT  277.475 0.17 277.735 10.48 ;
        RECT  277.985 0.17 278.245 10.99 ;
        RECT  276.48 118.025 276.68 118.755 ;
        RECT  277.3 118.025 277.5 118.755 ;
        RECT  278.495 0.17 279.265 0.94 ;
        RECT  278.495 0.17 278.755 8.7 ;
        RECT  279.005 0.17 279.265 12.9 ;
        RECT  277.795 118.025 277.995 118.755 ;
        RECT  278.295 118.025 278.495 118.755 ;
        RECT  278.795 118.025 278.995 118.755 ;
        RECT  279.29 118.025 279.49 118.755 ;
        RECT  279.515 0.52 279.775 2.485 ;
        RECT  280.11 118.025 280.31 118.755 ;
        RECT  280.38 0.52 280.64 14.11 ;
        RECT  280.605 118.025 280.805 118.755 ;
        RECT  280.89 0.52 281.15 2.335 ;
        RECT  281.105 118.025 281.305 118.755 ;
        RECT  281.605 118.025 281.805 118.755 ;
        RECT  282.1 118.025 282.3 118.755 ;
        RECT  284.29 0.52 284.55 5.16 ;
        RECT  283.77 4.9 284.55 5.16 ;
        RECT  283.77 4.9 284.03 6.64 ;
        RECT  282.92 118.025 283.12 118.755 ;
        RECT  283.415 118.025 283.615 118.755 ;
        RECT  283.915 118.025 284.115 118.755 ;
        RECT  284.415 118.025 284.615 118.755 ;
        RECT  284.91 118.025 285.11 118.755 ;
        RECT  285.655 0.17 286.425 0.94 ;
        RECT  285.655 0.17 285.915 12.9 ;
        RECT  286.165 0.17 286.425 12.9 ;
        RECT  285.145 0.52 285.405 5.815 ;
        RECT  285.73 118.025 285.93 118.755 ;
        RECT  286.675 0.17 287.445 0.43 ;
        RECT  286.675 0.17 286.935 11.5 ;
        RECT  287.185 0.17 287.445 11.5 ;
        RECT  286.225 118.025 286.425 118.755 ;
        RECT  286.725 118.025 286.925 118.755 ;
        RECT  287.225 118.025 287.425 118.755 ;
        RECT  288.715 0.17 289.485 0.43 ;
        RECT  288.715 0.17 288.975 10.48 ;
        RECT  289.225 0.17 289.485 10.99 ;
        RECT  287.72 118.025 287.92 118.755 ;
        RECT  288.54 118.025 288.74 118.755 ;
        RECT  289.735 0.17 290.505 0.94 ;
        RECT  289.735 0.17 289.995 8.7 ;
        RECT  290.245 0.17 290.505 12.9 ;
        RECT  289.035 118.025 289.235 118.755 ;
        RECT  289.535 118.025 289.735 118.755 ;
        RECT  290.035 118.025 290.235 118.755 ;
        RECT  290.53 118.025 290.73 118.755 ;
        RECT  290.755 0.52 291.015 2.485 ;
        RECT  291.35 118.025 291.55 118.755 ;
        RECT  291.62 0.52 291.88 14.11 ;
        RECT  291.845 118.025 292.045 118.755 ;
        RECT  292.13 0.52 292.39 2.335 ;
        RECT  292.345 118.025 292.545 118.755 ;
        RECT  292.845 118.025 293.045 118.755 ;
        RECT  293.34 118.025 293.54 118.755 ;
        RECT  295.53 0.52 295.79 5.16 ;
        RECT  295.01 4.9 295.79 5.16 ;
        RECT  295.01 4.9 295.27 6.64 ;
        RECT  294.16 118.025 294.36 118.755 ;
        RECT  294.655 118.025 294.855 118.755 ;
        RECT  295.155 118.025 295.355 118.755 ;
        RECT  295.655 118.025 295.855 118.755 ;
        RECT  296.15 118.025 296.35 118.755 ;
        RECT  296.895 0.17 297.665 0.94 ;
        RECT  296.895 0.17 297.155 12.9 ;
        RECT  297.405 0.17 297.665 12.9 ;
        RECT  296.385 0.52 296.645 5.815 ;
        RECT  296.97 118.025 297.17 118.755 ;
        RECT  297.915 0.17 298.685 0.43 ;
        RECT  297.915 0.17 298.175 11.5 ;
        RECT  298.425 0.17 298.685 11.5 ;
        RECT  297.465 118.025 297.665 118.755 ;
        RECT  297.965 118.025 298.165 118.755 ;
        RECT  298.465 118.025 298.665 118.755 ;
        RECT  299.955 0.17 300.725 0.43 ;
        RECT  299.955 0.17 300.215 10.48 ;
        RECT  300.465 0.17 300.725 10.99 ;
        RECT  298.96 118.025 299.16 118.755 ;
        RECT  299.78 118.025 299.98 118.755 ;
        RECT  300.975 0.17 301.745 0.94 ;
        RECT  300.975 0.17 301.235 8.7 ;
        RECT  301.485 0.17 301.745 12.9 ;
        RECT  300.275 118.025 300.475 118.755 ;
        RECT  300.775 118.025 300.975 118.755 ;
        RECT  301.275 118.025 301.475 118.755 ;
        RECT  301.77 118.025 301.97 118.755 ;
        RECT  301.995 0.52 302.255 2.485 ;
        RECT  302.59 118.025 302.79 118.755 ;
        RECT  302.86 0.52 303.12 14.11 ;
        RECT  303.085 118.025 303.285 118.755 ;
        RECT  303.37 0.52 303.63 2.335 ;
        RECT  303.585 118.025 303.785 118.755 ;
        RECT  304.085 118.025 304.285 118.755 ;
        RECT  304.58 118.025 304.78 118.755 ;
        RECT  306.77 0.52 307.03 5.16 ;
        RECT  306.25 4.9 307.03 5.16 ;
        RECT  306.25 4.9 306.51 6.64 ;
        RECT  305.4 118.025 305.6 118.755 ;
        RECT  305.895 118.025 306.095 118.755 ;
        RECT  306.395 118.025 306.595 118.755 ;
        RECT  306.895 118.025 307.095 118.755 ;
        RECT  307.39 118.025 307.59 118.755 ;
        RECT  308.135 0.17 308.905 0.94 ;
        RECT  308.135 0.17 308.395 12.9 ;
        RECT  308.645 0.17 308.905 12.9 ;
        RECT  307.625 0.52 307.885 5.815 ;
        RECT  308.21 118.025 308.41 118.755 ;
        RECT  309.155 0.17 309.925 0.43 ;
        RECT  309.155 0.17 309.415 11.5 ;
        RECT  309.665 0.17 309.925 11.5 ;
        RECT  308.705 118.025 308.905 118.755 ;
        RECT  309.205 118.025 309.405 118.755 ;
        RECT  309.705 118.025 309.905 118.755 ;
        RECT  311.195 0.17 311.965 0.43 ;
        RECT  311.195 0.17 311.455 10.48 ;
        RECT  311.705 0.17 311.965 10.99 ;
        RECT  310.2 118.025 310.4 118.755 ;
        RECT  311.02 118.025 311.22 118.755 ;
        RECT  312.215 0.17 312.985 0.94 ;
        RECT  312.215 0.17 312.475 8.7 ;
        RECT  312.725 0.17 312.985 12.9 ;
        RECT  311.515 118.025 311.715 118.755 ;
        RECT  312.015 118.025 312.215 118.755 ;
        RECT  312.515 118.025 312.715 118.755 ;
        RECT  313.01 118.025 313.21 118.755 ;
        RECT  313.235 0.52 313.495 2.485 ;
        RECT  313.83 118.025 314.03 118.755 ;
        RECT  314.1 0.52 314.36 14.11 ;
        RECT  314.325 118.025 314.525 118.755 ;
        RECT  314.61 0.52 314.87 2.335 ;
        RECT  314.825 118.025 315.025 118.755 ;
        RECT  315.325 118.025 315.525 118.755 ;
        RECT  315.82 118.025 316.02 118.755 ;
        RECT  318.01 0.52 318.27 5.16 ;
        RECT  317.49 4.9 318.27 5.16 ;
        RECT  317.49 4.9 317.75 6.64 ;
        RECT  316.64 118.025 316.84 118.755 ;
        RECT  317.135 118.025 317.335 118.755 ;
        RECT  317.635 118.025 317.835 118.755 ;
        RECT  318.135 118.025 318.335 118.755 ;
        RECT  318.63 118.025 318.83 118.755 ;
        RECT  319.375 0.17 320.145 0.94 ;
        RECT  319.375 0.17 319.635 12.9 ;
        RECT  319.885 0.17 320.145 12.9 ;
        RECT  318.865 0.52 319.125 5.815 ;
        RECT  319.45 118.025 319.65 118.755 ;
        RECT  320.395 0.17 321.165 0.43 ;
        RECT  320.395 0.17 320.655 11.5 ;
        RECT  320.905 0.17 321.165 11.5 ;
        RECT  319.945 118.025 320.145 118.755 ;
        RECT  320.445 118.025 320.645 118.755 ;
        RECT  320.945 118.025 321.145 118.755 ;
        RECT  322.435 0.17 323.205 0.43 ;
        RECT  322.435 0.17 322.695 10.48 ;
        RECT  322.945 0.17 323.205 10.99 ;
        RECT  321.44 118.025 321.64 118.755 ;
        RECT  322.26 118.025 322.46 118.755 ;
        RECT  323.455 0.17 324.225 0.94 ;
        RECT  323.455 0.17 323.715 8.7 ;
        RECT  323.965 0.17 324.225 12.9 ;
        RECT  322.755 118.025 322.955 118.755 ;
        RECT  323.255 118.025 323.455 118.755 ;
        RECT  323.755 118.025 323.955 118.755 ;
        RECT  324.25 118.025 324.45 118.755 ;
        RECT  324.475 0.52 324.735 2.485 ;
        RECT  325.07 118.025 325.27 118.755 ;
        RECT  325.34 0.52 325.6 14.11 ;
        RECT  325.565 118.025 325.765 118.755 ;
        RECT  325.85 0.52 326.11 2.335 ;
        RECT  326.065 118.025 326.265 118.755 ;
        RECT  326.565 118.025 326.765 118.755 ;
        RECT  327.06 118.025 327.26 118.755 ;
        RECT  329.25 0.52 329.51 5.16 ;
        RECT  328.73 4.9 329.51 5.16 ;
        RECT  328.73 4.9 328.99 6.64 ;
        RECT  327.88 118.025 328.08 118.755 ;
        RECT  328.375 118.025 328.575 118.755 ;
        RECT  328.875 118.025 329.075 118.755 ;
        RECT  329.375 118.025 329.575 118.755 ;
        RECT  329.87 118.025 330.07 118.755 ;
        RECT  330.615 0.17 331.385 0.94 ;
        RECT  330.615 0.17 330.875 12.9 ;
        RECT  331.125 0.17 331.385 12.9 ;
        RECT  330.105 0.52 330.365 5.815 ;
        RECT  330.69 118.025 330.89 118.755 ;
        RECT  331.635 0.17 332.405 0.43 ;
        RECT  331.635 0.17 331.895 11.5 ;
        RECT  332.145 0.17 332.405 11.5 ;
        RECT  331.185 118.025 331.385 118.755 ;
        RECT  331.685 118.025 331.885 118.755 ;
        RECT  332.185 118.025 332.385 118.755 ;
        RECT  333.675 0.17 334.445 0.43 ;
        RECT  333.675 0.17 333.935 10.48 ;
        RECT  334.185 0.17 334.445 10.99 ;
        RECT  332.68 118.025 332.88 118.755 ;
        RECT  333.5 118.025 333.7 118.755 ;
        RECT  334.695 0.17 335.465 0.94 ;
        RECT  334.695 0.17 334.955 8.7 ;
        RECT  335.205 0.17 335.465 12.9 ;
        RECT  333.995 118.025 334.195 118.755 ;
        RECT  334.495 118.025 334.695 118.755 ;
        RECT  334.995 118.025 335.195 118.755 ;
        RECT  335.49 118.025 335.69 118.755 ;
        RECT  335.715 0.52 335.975 2.485 ;
        RECT  336.31 118.025 336.51 118.755 ;
        RECT  336.58 0.52 336.84 14.11 ;
        RECT  336.805 118.025 337.005 118.755 ;
        RECT  337.09 0.52 337.35 2.335 ;
        RECT  337.305 118.025 337.505 118.755 ;
        RECT  337.805 118.025 338.005 118.755 ;
        RECT  338.3 118.025 338.5 118.755 ;
        RECT  340.49 0.52 340.75 5.16 ;
        RECT  339.97 4.9 340.75 5.16 ;
        RECT  339.97 4.9 340.23 6.64 ;
        RECT  339.12 118.025 339.32 118.755 ;
        RECT  339.615 118.025 339.815 118.755 ;
        RECT  340.115 118.025 340.315 118.755 ;
        RECT  340.615 118.025 340.815 118.755 ;
        RECT  341.11 118.025 341.31 118.755 ;
        RECT  341.855 0.17 342.625 0.94 ;
        RECT  341.855 0.17 342.115 12.9 ;
        RECT  342.365 0.17 342.625 12.9 ;
        RECT  341.345 0.52 341.605 5.815 ;
        RECT  341.93 118.025 342.13 118.755 ;
        RECT  342.875 0.17 343.645 0.43 ;
        RECT  342.875 0.17 343.135 11.5 ;
        RECT  343.385 0.17 343.645 11.5 ;
        RECT  342.425 118.025 342.625 118.755 ;
        RECT  342.925 118.025 343.125 118.755 ;
        RECT  343.425 118.025 343.625 118.755 ;
        RECT  344.915 0.17 345.685 0.43 ;
        RECT  344.915 0.17 345.175 10.48 ;
        RECT  345.425 0.17 345.685 10.99 ;
        RECT  343.92 118.025 344.12 118.755 ;
        RECT  344.74 118.025 344.94 118.755 ;
        RECT  345.935 0.17 346.705 0.94 ;
        RECT  345.935 0.17 346.195 8.7 ;
        RECT  346.445 0.17 346.705 12.9 ;
        RECT  345.235 118.025 345.435 118.755 ;
        RECT  345.735 118.025 345.935 118.755 ;
        RECT  346.235 118.025 346.435 118.755 ;
        RECT  346.73 118.025 346.93 118.755 ;
        RECT  346.955 0.52 347.215 2.485 ;
        RECT  347.55 118.025 347.75 118.755 ;
        RECT  347.82 0.52 348.08 14.11 ;
        RECT  348.045 118.025 348.245 118.755 ;
        RECT  348.33 0.52 348.59 2.335 ;
        RECT  348.545 118.025 348.745 118.755 ;
        RECT  349.045 118.025 349.245 118.755 ;
        RECT  349.54 118.025 349.74 118.755 ;
        RECT  351.73 0.52 351.99 5.16 ;
        RECT  351.21 4.9 351.99 5.16 ;
        RECT  351.21 4.9 351.47 6.64 ;
        RECT  350.36 118.025 350.56 118.755 ;
        RECT  350.855 118.025 351.055 118.755 ;
        RECT  351.355 118.025 351.555 118.755 ;
        RECT  351.855 118.025 352.055 118.755 ;
        RECT  352.35 118.025 352.55 118.755 ;
        RECT  353.095 0.17 353.865 0.94 ;
        RECT  353.095 0.17 353.355 12.9 ;
        RECT  353.605 0.17 353.865 12.9 ;
        RECT  352.585 0.52 352.845 5.815 ;
        RECT  353.17 118.025 353.37 118.755 ;
        RECT  354.115 0.17 354.885 0.43 ;
        RECT  354.115 0.17 354.375 11.5 ;
        RECT  354.625 0.17 354.885 11.5 ;
        RECT  353.665 118.025 353.865 118.755 ;
        RECT  354.165 118.025 354.365 118.755 ;
        RECT  354.665 118.025 354.865 118.755 ;
        RECT  356.155 0.17 356.925 0.43 ;
        RECT  356.155 0.17 356.415 10.48 ;
        RECT  356.665 0.17 356.925 10.99 ;
        RECT  355.16 118.025 355.36 118.755 ;
        RECT  355.98 118.025 356.18 118.755 ;
        RECT  357.175 0.17 357.945 0.94 ;
        RECT  357.175 0.17 357.435 8.7 ;
        RECT  357.685 0.17 357.945 12.9 ;
        RECT  356.475 118.025 356.675 118.755 ;
        RECT  356.975 118.025 357.175 118.755 ;
        RECT  357.475 118.025 357.675 118.755 ;
        RECT  357.97 118.025 358.17 118.755 ;
        RECT  358.195 0.52 358.455 2.485 ;
        RECT  358.79 118.025 358.99 118.755 ;
        RECT  359.06 0.52 359.32 14.11 ;
        RECT  359.285 118.025 359.485 118.755 ;
        RECT  359.57 0.52 359.83 2.335 ;
        RECT  359.785 118.025 359.985 118.755 ;
        RECT  360.285 118.025 360.485 118.755 ;
        RECT  362.275 0.17 363.045 0.43 ;
        RECT  362.275 0.17 362.535 8.7 ;
        RECT  362.785 0.17 363.045 8.7 ;
        RECT  363.295 0.17 364.065 0.94 ;
        RECT  363.295 0.17 363.555 8.7 ;
        RECT  363.805 0.17 364.065 8.7 ;
        RECT  364.315 0.17 365.085 0.43 ;
        RECT  364.315 0.17 364.575 8.7 ;
        RECT  364.825 0.17 365.085 8.7 ;
        RECT  365.335 0.17 366.105 0.94 ;
        RECT  365.335 0.17 365.595 8.7 ;
        RECT  365.845 0.17 366.105 8.7 ;
        RECT  366.355 0.17 367.125 0.43 ;
        RECT  366.355 0.17 366.615 8.7 ;
        RECT  366.865 0.17 367.125 8.7 ;
        RECT  367.375 0.17 368.145 0.94 ;
        RECT  367.375 0.17 367.635 8.7 ;
        RECT  367.885 0.17 368.145 8.7 ;
        RECT  368.395 0.17 369.165 0.43 ;
        RECT  368.395 0.17 368.655 8.7 ;
        RECT  368.905 0.17 369.165 8.7 ;
        RECT  369.415 0.17 370.185 0.94 ;
        RECT  369.415 0.17 369.675 8.7 ;
        RECT  369.925 0.17 370.185 8.7 ;
        RECT  370.435 0.17 371.205 0.43 ;
        RECT  370.435 0.17 370.695 8.7 ;
        RECT  370.945 0.17 371.205 8.7 ;
        RECT  371.455 0.17 372.225 0.94 ;
        RECT  371.455 0.17 371.715 8.7 ;
        RECT  371.965 0.17 372.225 8.7 ;
        RECT  360.78 118.025 360.98 118.755 ;
        RECT  361.6 118.025 361.8 118.755 ;
        RECT  362.595 118.025 362.795 118.755 ;
        RECT  374.16 0.17 374.93 0.94 ;
        RECT  374.16 0.17 374.42 8.7 ;
        RECT  374.67 0.17 374.93 8.7 ;
        RECT  372.63 0.3 372.89 8.7 ;
        RECT  373.14 0 373.4 8.7 ;
        RECT  373.65 0 373.91 8.7 ;
        RECT  375.18 0 375.44 8.7 ;
        RECT  375.69 0 375.95 8.7 ;
        RECT  376.2 0.52 376.46 8.7 ;
        RECT  376.71 0.52 376.97 8.7 ;
        RECT  377.22 0.52 377.48 8.7 ;
        RECT  379.26 0.17 380.03 0.94 ;
        RECT  379.26 0.17 379.52 8.7 ;
        RECT  379.77 0.17 380.03 8.7 ;
        RECT  380.28 0.17 381.05 0.43 ;
        RECT  380.28 0.17 380.54 8.7 ;
        RECT  380.79 0.17 381.05 8.7 ;
        RECT  377.73 0.52 377.99 8.7 ;
        RECT  378.24 0 378.5 8.7 ;
        RECT  378.75 0 379.01 8.7 ;
        RECT  381.3 0.3 381.56 8.7 ;
        RECT  381.81 0.3 382.07 8.7 ;
        RECT  383.85 0.17 384.62 0.94 ;
        RECT  383.85 0.17 384.11 8.7 ;
        RECT  384.36 0.17 384.62 8.7 ;
        RECT  382.32 0.3 382.58 8.7 ;
        RECT  382.83 0.3 383.09 8.7 ;
        RECT  383.34 0.3 383.6 8.7 ;
        RECT  384.87 0.52 385.13 8.7 ;
        RECT  385.38 0.52 385.64 8.7 ;
        RECT  385.89 0.3 386.15 8.7 ;
        RECT  386.4 0.52 386.66 8.7 ;
        RECT  386.91 0.52 387.17 8.7 ;
        RECT  387.42 0.3 387.68 8.7 ;
        RECT  387.93 0.52 388.19 8.7 ;
        RECT  388.44 0.52 388.7 8.7 ;
        RECT  388.95 0.52 389.21 8.7 ;
        RECT  389.46 0.52 389.72 8.7 ;
        RECT  389.97 0.52 390.23 8.7 ;
        RECT  390.48 0.3 390.74 8.7 ;
        RECT  390.99 0.52 391.25 8.7 ;
        RECT  391.5 0.52 391.76 8.7 ;
        RECT  392.01 0.3 392.27 8.7 ;
        RECT  394.05 0.17 394.82 0.94 ;
        RECT  394.05 0.17 394.31 8.7 ;
        RECT  394.56 0.17 394.82 8.7 ;
        RECT  392.52 0.52 392.78 8.7 ;
        RECT  393.03 0.52 393.29 8.7 ;
        RECT  393.54 0.3 393.8 8.7 ;
        RECT  395.07 0.52 395.33 8.7 ;
        RECT  395.58 0.52 395.84 8.7 ;
        RECT  396.09 0.52 396.35 8.7 ;
        RECT  396.6 0.52 396.86 8.7 ;
        RECT  397.11 0.52 397.37 8.7 ;
        RECT  397.62 0.52 397.88 8.7 ;
        RECT  398.13 0.52 398.39 8.7 ;
        RECT  400.17 0.17 400.94 0.94 ;
        RECT  400.17 0.17 400.43 8.7 ;
        RECT  400.68 0.17 400.94 8.7 ;
        RECT  398.64 0.52 398.9 8.7 ;
        RECT  399.15 0 399.41 8.7 ;
        RECT  399.66 0 399.92 8.7 ;
        RECT  401.19 0 401.45 8.7 ;
        RECT  403.23 0.17 404 0.43 ;
        RECT  403.23 0.17 403.49 8.7 ;
        RECT  403.74 0.17 404 8.7 ;
        RECT  401.7 0 401.96 8.7 ;
        RECT  402.21 0.3 402.47 8.7 ;
        RECT  402.72 0.3 402.98 8.7 ;
        RECT  404.25 0.3 404.51 8.7 ;
        RECT  404.76 0.3 405.02 8.7 ;
        RECT  405.27 0.3 405.53 8.7 ;
        RECT  405.78 0.3 406.04 8.7 ;
        RECT  406.29 0 406.55 8.7 ;
        RECT  406.8 0 407.06 8.7 ;
        RECT  408.84 0.17 409.61 0.43 ;
        RECT  408.84 0.17 409.1 8.7 ;
        RECT  409.35 0.17 409.61 8.7 ;
        RECT  409.86 0.17 410.63 0.94 ;
        RECT  409.86 0.17 410.12 25.5 ;
        RECT  410.37 0.17 410.63 33.9 ;
        RECT  410.88 0.17 411.65 0.43 ;
        RECT  410.88 0.17 411.14 8.7 ;
        RECT  411.39 0.17 411.65 8.7 ;
        RECT  412.255 0.17 413.025 0.94 ;
        RECT  412.255 0.17 412.515 8.7 ;
        RECT  412.765 0.17 413.025 8.7 ;
        RECT  413.275 0.17 414.045 0.43 ;
        RECT  413.275 0.17 413.535 8.7 ;
        RECT  413.785 0.17 414.045 8.7 ;
        RECT  414.295 0.17 415.065 0.94 ;
        RECT  414.295 0.17 414.555 8.7 ;
        RECT  414.805 0.17 415.065 8.7 ;
        RECT  415.315 0.17 416.085 0.43 ;
        RECT  415.315 0.17 415.575 8.7 ;
        RECT  415.825 0.17 416.085 8.7 ;
        RECT  416.335 0.17 417.105 0.94 ;
        RECT  416.335 0.17 416.595 8.7 ;
        RECT  416.845 0.17 417.105 8.7 ;
        RECT  417.355 0.17 418.125 0.43 ;
        RECT  417.355 0.17 417.615 8.7 ;
        RECT  417.865 0.17 418.125 8.7 ;
        RECT  418.375 0.17 419.145 0.94 ;
        RECT  418.375 0.17 418.635 8.7 ;
        RECT  418.885 0.17 419.145 8.7 ;
        RECT  419.395 0.17 420.165 0.43 ;
        RECT  419.395 0.17 419.655 8.7 ;
        RECT  419.905 0.17 420.165 8.7 ;
        RECT  420.415 0.17 421.185 0.94 ;
        RECT  420.415 0.17 420.675 8.7 ;
        RECT  420.925 0.17 421.185 8.7 ;
        RECT  407.31 0.3 407.57 8.7 ;
        RECT  421.435 0.17 422.205 0.43 ;
        RECT  421.435 0.17 421.695 8.7 ;
        RECT  421.945 0.17 422.205 8.7 ;
        RECT  407.82 0.3 408.08 8.7 ;
        RECT  408.33 0.52 408.59 8.7 ;
        RECT  421.685 118.025 421.885 118.755 ;
        RECT  422.68 118.025 422.88 118.755 ;
        RECT  423.5 118.025 423.7 118.755 ;
        RECT  423.995 118.025 424.195 118.755 ;
        RECT  424.495 118.025 424.695 118.755 ;
        RECT  424.65 0.52 424.91 2.335 ;
        RECT  424.995 118.025 425.195 118.755 ;
        RECT  425.16 0.52 425.42 14.11 ;
        RECT  425.49 118.025 425.69 118.755 ;
        RECT  426.535 0.17 427.305 0.94 ;
        RECT  427.045 0.17 427.305 8.7 ;
        RECT  426.535 0.17 426.795 12.9 ;
        RECT  426.025 0.52 426.285 2.485 ;
        RECT  426.31 118.025 426.51 118.755 ;
        RECT  427.555 0.17 428.325 0.43 ;
        RECT  428.065 0.17 428.325 10.48 ;
        RECT  427.555 0.17 427.815 10.99 ;
        RECT  426.805 118.025 427.005 118.755 ;
        RECT  427.305 118.025 427.505 118.755 ;
        RECT  427.805 118.025 428.005 118.755 ;
        RECT  428.3 118.025 428.5 118.755 ;
        RECT  429.595 0.17 430.365 0.43 ;
        RECT  429.595 0.17 429.855 11.5 ;
        RECT  430.105 0.17 430.365 11.5 ;
        RECT  429.12 118.025 429.32 118.755 ;
        RECT  429.615 118.025 429.815 118.755 ;
        RECT  430.615 0.17 431.385 0.94 ;
        RECT  430.615 0.17 430.875 12.9 ;
        RECT  431.125 0.17 431.385 12.9 ;
        RECT  430.115 118.025 430.315 118.755 ;
        RECT  430.615 118.025 430.815 118.755 ;
        RECT  431.11 118.025 431.31 118.755 ;
        RECT  431.635 0.52 431.895 5.815 ;
        RECT  432.49 0.52 432.75 5.16 ;
        RECT  432.49 4.9 433.27 5.16 ;
        RECT  433.01 4.9 433.27 6.64 ;
        RECT  431.93 118.025 432.13 118.755 ;
        RECT  432.425 118.025 432.625 118.755 ;
        RECT  432.925 118.025 433.125 118.755 ;
        RECT  433.425 118.025 433.625 118.755 ;
        RECT  433.92 118.025 434.12 118.755 ;
        RECT  434.74 118.025 434.94 118.755 ;
        RECT  435.235 118.025 435.435 118.755 ;
        RECT  435.735 118.025 435.935 118.755 ;
        RECT  435.89 0.52 436.15 2.335 ;
        RECT  436.235 118.025 436.435 118.755 ;
        RECT  436.4 0.52 436.66 14.11 ;
        RECT  436.73 118.025 436.93 118.755 ;
        RECT  437.775 0.17 438.545 0.94 ;
        RECT  438.285 0.17 438.545 8.7 ;
        RECT  437.775 0.17 438.035 12.9 ;
        RECT  437.265 0.52 437.525 2.485 ;
        RECT  437.55 118.025 437.75 118.755 ;
        RECT  438.795 0.17 439.565 0.43 ;
        RECT  439.305 0.17 439.565 10.48 ;
        RECT  438.795 0.17 439.055 10.99 ;
        RECT  438.045 118.025 438.245 118.755 ;
        RECT  438.545 118.025 438.745 118.755 ;
        RECT  439.045 118.025 439.245 118.755 ;
        RECT  439.54 118.025 439.74 118.755 ;
        RECT  440.835 0.17 441.605 0.43 ;
        RECT  440.835 0.17 441.095 11.5 ;
        RECT  441.345 0.17 441.605 11.5 ;
        RECT  440.36 118.025 440.56 118.755 ;
        RECT  440.855 118.025 441.055 118.755 ;
        RECT  441.855 0.17 442.625 0.94 ;
        RECT  441.855 0.17 442.115 12.9 ;
        RECT  442.365 0.17 442.625 12.9 ;
        RECT  441.355 118.025 441.555 118.755 ;
        RECT  441.855 118.025 442.055 118.755 ;
        RECT  442.35 118.025 442.55 118.755 ;
        RECT  442.875 0.52 443.135 5.815 ;
        RECT  443.73 0.52 443.99 5.16 ;
        RECT  443.73 4.9 444.51 5.16 ;
        RECT  444.25 4.9 444.51 6.64 ;
        RECT  443.17 118.025 443.37 118.755 ;
        RECT  443.665 118.025 443.865 118.755 ;
        RECT  444.165 118.025 444.365 118.755 ;
        RECT  444.665 118.025 444.865 118.755 ;
        RECT  445.16 118.025 445.36 118.755 ;
        RECT  445.98 118.025 446.18 118.755 ;
        RECT  446.475 118.025 446.675 118.755 ;
        RECT  446.975 118.025 447.175 118.755 ;
        RECT  447.13 0.52 447.39 2.335 ;
        RECT  447.475 118.025 447.675 118.755 ;
        RECT  447.64 0.52 447.9 14.11 ;
        RECT  447.97 118.025 448.17 118.755 ;
        RECT  449.015 0.17 449.785 0.94 ;
        RECT  449.525 0.17 449.785 8.7 ;
        RECT  449.015 0.17 449.275 12.9 ;
        RECT  448.505 0.52 448.765 2.485 ;
        RECT  448.79 118.025 448.99 118.755 ;
        RECT  450.035 0.17 450.805 0.43 ;
        RECT  450.545 0.17 450.805 10.48 ;
        RECT  450.035 0.17 450.295 10.99 ;
        RECT  449.285 118.025 449.485 118.755 ;
        RECT  449.785 118.025 449.985 118.755 ;
        RECT  450.285 118.025 450.485 118.755 ;
        RECT  450.78 118.025 450.98 118.755 ;
        RECT  452.075 0.17 452.845 0.43 ;
        RECT  452.075 0.17 452.335 11.5 ;
        RECT  452.585 0.17 452.845 11.5 ;
        RECT  451.6 118.025 451.8 118.755 ;
        RECT  452.095 118.025 452.295 118.755 ;
        RECT  453.095 0.17 453.865 0.94 ;
        RECT  453.095 0.17 453.355 12.9 ;
        RECT  453.605 0.17 453.865 12.9 ;
        RECT  452.595 118.025 452.795 118.755 ;
        RECT  453.095 118.025 453.295 118.755 ;
        RECT  453.59 118.025 453.79 118.755 ;
        RECT  454.115 0.52 454.375 5.815 ;
        RECT  454.97 0.52 455.23 5.16 ;
        RECT  454.97 4.9 455.75 5.16 ;
        RECT  455.49 4.9 455.75 6.64 ;
        RECT  454.41 118.025 454.61 118.755 ;
        RECT  454.905 118.025 455.105 118.755 ;
        RECT  455.405 118.025 455.605 118.755 ;
        RECT  455.905 118.025 456.105 118.755 ;
        RECT  456.4 118.025 456.6 118.755 ;
        RECT  457.22 118.025 457.42 118.755 ;
        RECT  457.715 118.025 457.915 118.755 ;
        RECT  458.215 118.025 458.415 118.755 ;
        RECT  458.37 0.52 458.63 2.335 ;
        RECT  458.715 118.025 458.915 118.755 ;
        RECT  458.88 0.52 459.14 14.11 ;
        RECT  459.21 118.025 459.41 118.755 ;
        RECT  460.255 0.17 461.025 0.94 ;
        RECT  460.765 0.17 461.025 8.7 ;
        RECT  460.255 0.17 460.515 12.9 ;
        RECT  459.745 0.52 460.005 2.485 ;
        RECT  460.03 118.025 460.23 118.755 ;
        RECT  461.275 0.17 462.045 0.43 ;
        RECT  461.785 0.17 462.045 10.48 ;
        RECT  461.275 0.17 461.535 10.99 ;
        RECT  460.525 118.025 460.725 118.755 ;
        RECT  461.025 118.025 461.225 118.755 ;
        RECT  461.525 118.025 461.725 118.755 ;
        RECT  462.02 118.025 462.22 118.755 ;
        RECT  463.315 0.17 464.085 0.43 ;
        RECT  463.315 0.17 463.575 11.5 ;
        RECT  463.825 0.17 464.085 11.5 ;
        RECT  462.84 118.025 463.04 118.755 ;
        RECT  463.335 118.025 463.535 118.755 ;
        RECT  464.335 0.17 465.105 0.94 ;
        RECT  464.335 0.17 464.595 12.9 ;
        RECT  464.845 0.17 465.105 12.9 ;
        RECT  463.835 118.025 464.035 118.755 ;
        RECT  464.335 118.025 464.535 118.755 ;
        RECT  464.83 118.025 465.03 118.755 ;
        RECT  465.355 0.52 465.615 5.815 ;
        RECT  466.21 0.52 466.47 5.16 ;
        RECT  466.21 4.9 466.99 5.16 ;
        RECT  466.73 4.9 466.99 6.64 ;
        RECT  465.65 118.025 465.85 118.755 ;
        RECT  466.145 118.025 466.345 118.755 ;
        RECT  466.645 118.025 466.845 118.755 ;
        RECT  467.145 118.025 467.345 118.755 ;
        RECT  467.64 118.025 467.84 118.755 ;
        RECT  468.46 118.025 468.66 118.755 ;
        RECT  468.955 118.025 469.155 118.755 ;
        RECT  469.455 118.025 469.655 118.755 ;
        RECT  469.61 0.52 469.87 2.335 ;
        RECT  469.955 118.025 470.155 118.755 ;
        RECT  470.12 0.52 470.38 14.11 ;
        RECT  470.45 118.025 470.65 118.755 ;
        RECT  471.495 0.17 472.265 0.94 ;
        RECT  472.005 0.17 472.265 8.7 ;
        RECT  471.495 0.17 471.755 12.9 ;
        RECT  470.985 0.52 471.245 2.485 ;
        RECT  471.27 118.025 471.47 118.755 ;
        RECT  472.515 0.17 473.285 0.43 ;
        RECT  473.025 0.17 473.285 10.48 ;
        RECT  472.515 0.17 472.775 10.99 ;
        RECT  471.765 118.025 471.965 118.755 ;
        RECT  472.265 118.025 472.465 118.755 ;
        RECT  472.765 118.025 472.965 118.755 ;
        RECT  473.26 118.025 473.46 118.755 ;
        RECT  474.555 0.17 475.325 0.43 ;
        RECT  474.555 0.17 474.815 11.5 ;
        RECT  475.065 0.17 475.325 11.5 ;
        RECT  474.08 118.025 474.28 118.755 ;
        RECT  474.575 118.025 474.775 118.755 ;
        RECT  475.575 0.17 476.345 0.94 ;
        RECT  475.575 0.17 475.835 12.9 ;
        RECT  476.085 0.17 476.345 12.9 ;
        RECT  475.075 118.025 475.275 118.755 ;
        RECT  475.575 118.025 475.775 118.755 ;
        RECT  476.07 118.025 476.27 118.755 ;
        RECT  476.595 0.52 476.855 5.815 ;
        RECT  477.45 0.52 477.71 5.16 ;
        RECT  477.45 4.9 478.23 5.16 ;
        RECT  477.97 4.9 478.23 6.64 ;
        RECT  476.89 118.025 477.09 118.755 ;
        RECT  477.385 118.025 477.585 118.755 ;
        RECT  477.885 118.025 478.085 118.755 ;
        RECT  478.385 118.025 478.585 118.755 ;
        RECT  478.88 118.025 479.08 118.755 ;
        RECT  479.7 118.025 479.9 118.755 ;
        RECT  480.195 118.025 480.395 118.755 ;
        RECT  480.695 118.025 480.895 118.755 ;
        RECT  480.85 0.52 481.11 2.335 ;
        RECT  481.195 118.025 481.395 118.755 ;
        RECT  481.36 0.52 481.62 14.11 ;
        RECT  481.69 118.025 481.89 118.755 ;
        RECT  482.735 0.17 483.505 0.94 ;
        RECT  483.245 0.17 483.505 8.7 ;
        RECT  482.735 0.17 482.995 12.9 ;
        RECT  482.225 0.52 482.485 2.485 ;
        RECT  482.51 118.025 482.71 118.755 ;
        RECT  483.755 0.17 484.525 0.43 ;
        RECT  484.265 0.17 484.525 10.48 ;
        RECT  483.755 0.17 484.015 10.99 ;
        RECT  483.005 118.025 483.205 118.755 ;
        RECT  483.505 118.025 483.705 118.755 ;
        RECT  484.005 118.025 484.205 118.755 ;
        RECT  484.5 118.025 484.7 118.755 ;
        RECT  485.795 0.17 486.565 0.43 ;
        RECT  485.795 0.17 486.055 11.5 ;
        RECT  486.305 0.17 486.565 11.5 ;
        RECT  485.32 118.025 485.52 118.755 ;
        RECT  485.815 118.025 486.015 118.755 ;
        RECT  486.815 0.17 487.585 0.94 ;
        RECT  486.815 0.17 487.075 12.9 ;
        RECT  487.325 0.17 487.585 12.9 ;
        RECT  486.315 118.025 486.515 118.755 ;
        RECT  486.815 118.025 487.015 118.755 ;
        RECT  487.31 118.025 487.51 118.755 ;
        RECT  487.835 0.52 488.095 5.815 ;
        RECT  488.69 0.52 488.95 5.16 ;
        RECT  488.69 4.9 489.47 5.16 ;
        RECT  489.21 4.9 489.47 6.64 ;
        RECT  488.13 118.025 488.33 118.755 ;
        RECT  488.625 118.025 488.825 118.755 ;
        RECT  489.125 118.025 489.325 118.755 ;
        RECT  489.625 118.025 489.825 118.755 ;
        RECT  490.12 118.025 490.32 118.755 ;
        RECT  490.94 118.025 491.14 118.755 ;
        RECT  491.435 118.025 491.635 118.755 ;
        RECT  491.935 118.025 492.135 118.755 ;
        RECT  492.09 0.52 492.35 2.335 ;
        RECT  492.435 118.025 492.635 118.755 ;
        RECT  492.6 0.52 492.86 14.11 ;
        RECT  492.93 118.025 493.13 118.755 ;
        RECT  493.975 0.17 494.745 0.94 ;
        RECT  494.485 0.17 494.745 8.7 ;
        RECT  493.975 0.17 494.235 12.9 ;
        RECT  493.465 0.52 493.725 2.485 ;
        RECT  493.75 118.025 493.95 118.755 ;
        RECT  494.995 0.17 495.765 0.43 ;
        RECT  495.505 0.17 495.765 10.48 ;
        RECT  494.995 0.17 495.255 10.99 ;
        RECT  494.245 118.025 494.445 118.755 ;
        RECT  494.745 118.025 494.945 118.755 ;
        RECT  495.245 118.025 495.445 118.755 ;
        RECT  495.74 118.025 495.94 118.755 ;
        RECT  497.035 0.17 497.805 0.43 ;
        RECT  497.035 0.17 497.295 11.5 ;
        RECT  497.545 0.17 497.805 11.5 ;
        RECT  496.56 118.025 496.76 118.755 ;
        RECT  497.055 118.025 497.255 118.755 ;
        RECT  498.055 0.17 498.825 0.94 ;
        RECT  498.055 0.17 498.315 12.9 ;
        RECT  498.565 0.17 498.825 12.9 ;
        RECT  497.555 118.025 497.755 118.755 ;
        RECT  498.055 118.025 498.255 118.755 ;
        RECT  498.55 118.025 498.75 118.755 ;
        RECT  499.075 0.52 499.335 5.815 ;
        RECT  499.93 0.52 500.19 5.16 ;
        RECT  499.93 4.9 500.71 5.16 ;
        RECT  500.45 4.9 500.71 6.64 ;
        RECT  499.37 118.025 499.57 118.755 ;
        RECT  499.865 118.025 500.065 118.755 ;
        RECT  500.365 118.025 500.565 118.755 ;
        RECT  500.865 118.025 501.065 118.755 ;
        RECT  501.36 118.025 501.56 118.755 ;
        RECT  502.18 118.025 502.38 118.755 ;
        RECT  502.675 118.025 502.875 118.755 ;
        RECT  503.175 118.025 503.375 118.755 ;
        RECT  503.33 0.52 503.59 2.335 ;
        RECT  503.675 118.025 503.875 118.755 ;
        RECT  503.84 0.52 504.1 14.11 ;
        RECT  504.17 118.025 504.37 118.755 ;
        RECT  505.215 0.17 505.985 0.94 ;
        RECT  505.725 0.17 505.985 8.7 ;
        RECT  505.215 0.17 505.475 12.9 ;
        RECT  504.705 0.52 504.965 2.485 ;
        RECT  504.99 118.025 505.19 118.755 ;
        RECT  506.235 0.17 507.005 0.43 ;
        RECT  506.745 0.17 507.005 10.48 ;
        RECT  506.235 0.17 506.495 10.99 ;
        RECT  505.485 118.025 505.685 118.755 ;
        RECT  505.985 118.025 506.185 118.755 ;
        RECT  506.485 118.025 506.685 118.755 ;
        RECT  506.98 118.025 507.18 118.755 ;
        RECT  508.275 0.17 509.045 0.43 ;
        RECT  508.275 0.17 508.535 11.5 ;
        RECT  508.785 0.17 509.045 11.5 ;
        RECT  507.8 118.025 508 118.755 ;
        RECT  508.295 118.025 508.495 118.755 ;
        RECT  509.295 0.17 510.065 0.94 ;
        RECT  509.295 0.17 509.555 12.9 ;
        RECT  509.805 0.17 510.065 12.9 ;
        RECT  508.795 118.025 508.995 118.755 ;
        RECT  509.295 118.025 509.495 118.755 ;
        RECT  509.79 118.025 509.99 118.755 ;
        RECT  510.315 0.52 510.575 5.815 ;
        RECT  511.17 0.52 511.43 5.16 ;
        RECT  511.17 4.9 511.95 5.16 ;
        RECT  511.69 4.9 511.95 6.64 ;
        RECT  510.61 118.025 510.81 118.755 ;
        RECT  511.105 118.025 511.305 118.755 ;
        RECT  511.605 118.025 511.805 118.755 ;
        RECT  512.105 118.025 512.305 118.755 ;
        RECT  512.6 118.025 512.8 118.755 ;
        RECT  513.42 118.025 513.62 118.755 ;
        RECT  513.915 118.025 514.115 118.755 ;
        RECT  514.415 118.025 514.615 118.755 ;
        RECT  514.57 0.52 514.83 2.335 ;
        RECT  514.915 118.025 515.115 118.755 ;
        RECT  515.08 0.52 515.34 14.11 ;
        RECT  515.41 118.025 515.61 118.755 ;
        RECT  516.455 0.17 517.225 0.94 ;
        RECT  516.965 0.17 517.225 8.7 ;
        RECT  516.455 0.17 516.715 12.9 ;
        RECT  515.945 0.52 516.205 2.485 ;
        RECT  516.23 118.025 516.43 118.755 ;
        RECT  517.475 0.17 518.245 0.43 ;
        RECT  517.985 0.17 518.245 10.48 ;
        RECT  517.475 0.17 517.735 10.99 ;
        RECT  516.725 118.025 516.925 118.755 ;
        RECT  517.225 118.025 517.425 118.755 ;
        RECT  517.725 118.025 517.925 118.755 ;
        RECT  518.22 118.025 518.42 118.755 ;
        RECT  519.515 0.17 520.285 0.43 ;
        RECT  519.515 0.17 519.775 11.5 ;
        RECT  520.025 0.17 520.285 11.5 ;
        RECT  519.04 118.025 519.24 118.755 ;
        RECT  519.535 118.025 519.735 118.755 ;
        RECT  520.535 0.17 521.305 0.94 ;
        RECT  520.535 0.17 520.795 12.9 ;
        RECT  521.045 0.17 521.305 12.9 ;
        RECT  520.035 118.025 520.235 118.755 ;
        RECT  520.535 118.025 520.735 118.755 ;
        RECT  521.03 118.025 521.23 118.755 ;
        RECT  521.555 0.52 521.815 5.815 ;
        RECT  522.41 0.52 522.67 5.16 ;
        RECT  522.41 4.9 523.19 5.16 ;
        RECT  522.93 4.9 523.19 6.64 ;
        RECT  521.85 118.025 522.05 118.755 ;
        RECT  522.345 118.025 522.545 118.755 ;
        RECT  522.845 118.025 523.045 118.755 ;
        RECT  523.345 118.025 523.545 118.755 ;
        RECT  523.84 118.025 524.04 118.755 ;
        RECT  524.66 118.025 524.86 118.755 ;
        RECT  525.155 118.025 525.355 118.755 ;
        RECT  525.655 118.025 525.855 118.755 ;
        RECT  525.81 0.52 526.07 2.335 ;
        RECT  526.155 118.025 526.355 118.755 ;
        RECT  526.32 0.52 526.58 14.11 ;
        RECT  526.65 118.025 526.85 118.755 ;
        RECT  527.695 0.17 528.465 0.94 ;
        RECT  528.205 0.17 528.465 8.7 ;
        RECT  527.695 0.17 527.955 12.9 ;
        RECT  527.185 0.52 527.445 2.485 ;
        RECT  527.47 118.025 527.67 118.755 ;
        RECT  528.715 0.17 529.485 0.43 ;
        RECT  529.225 0.17 529.485 10.48 ;
        RECT  528.715 0.17 528.975 10.99 ;
        RECT  527.965 118.025 528.165 118.755 ;
        RECT  528.465 118.025 528.665 118.755 ;
        RECT  528.965 118.025 529.165 118.755 ;
        RECT  529.46 118.025 529.66 118.755 ;
        RECT  530.755 0.17 531.525 0.43 ;
        RECT  530.755 0.17 531.015 11.5 ;
        RECT  531.265 0.17 531.525 11.5 ;
        RECT  530.28 118.025 530.48 118.755 ;
        RECT  530.775 118.025 530.975 118.755 ;
        RECT  531.775 0.17 532.545 0.94 ;
        RECT  531.775 0.17 532.035 12.9 ;
        RECT  532.285 0.17 532.545 12.9 ;
        RECT  531.275 118.025 531.475 118.755 ;
        RECT  531.775 118.025 531.975 118.755 ;
        RECT  532.27 118.025 532.47 118.755 ;
        RECT  532.795 0.52 533.055 5.815 ;
        RECT  533.65 0.52 533.91 5.16 ;
        RECT  533.65 4.9 534.43 5.16 ;
        RECT  534.17 4.9 534.43 6.64 ;
        RECT  533.09 118.025 533.29 118.755 ;
        RECT  533.585 118.025 533.785 118.755 ;
        RECT  534.085 118.025 534.285 118.755 ;
        RECT  534.585 118.025 534.785 118.755 ;
        RECT  535.08 118.025 535.28 118.755 ;
        RECT  535.9 118.025 536.1 118.755 ;
        RECT  536.395 118.025 536.595 118.755 ;
        RECT  536.895 118.025 537.095 118.755 ;
        RECT  537.05 0.52 537.31 2.335 ;
        RECT  537.395 118.025 537.595 118.755 ;
        RECT  537.56 0.52 537.82 14.11 ;
        RECT  537.89 118.025 538.09 118.755 ;
        RECT  538.935 0.17 539.705 0.94 ;
        RECT  539.445 0.17 539.705 8.7 ;
        RECT  538.935 0.17 539.195 12.9 ;
        RECT  538.425 0.52 538.685 2.485 ;
        RECT  538.71 118.025 538.91 118.755 ;
        RECT  539.955 0.17 540.725 0.43 ;
        RECT  540.465 0.17 540.725 10.48 ;
        RECT  539.955 0.17 540.215 10.99 ;
        RECT  539.205 118.025 539.405 118.755 ;
        RECT  539.705 118.025 539.905 118.755 ;
        RECT  540.205 118.025 540.405 118.755 ;
        RECT  540.7 118.025 540.9 118.755 ;
        RECT  541.995 0.17 542.765 0.43 ;
        RECT  541.995 0.17 542.255 11.5 ;
        RECT  542.505 0.17 542.765 11.5 ;
        RECT  541.52 118.025 541.72 118.755 ;
        RECT  542.015 118.025 542.215 118.755 ;
        RECT  543.015 0.17 543.785 0.94 ;
        RECT  543.015 0.17 543.275 12.9 ;
        RECT  543.525 0.17 543.785 12.9 ;
        RECT  542.515 118.025 542.715 118.755 ;
        RECT  543.015 118.025 543.215 118.755 ;
        RECT  543.51 118.025 543.71 118.755 ;
        RECT  544.035 0.52 544.295 5.815 ;
        RECT  544.89 0.52 545.15 5.16 ;
        RECT  544.89 4.9 545.67 5.16 ;
        RECT  545.41 4.9 545.67 6.64 ;
        RECT  544.33 118.025 544.53 118.755 ;
        RECT  544.825 118.025 545.025 118.755 ;
        RECT  545.325 118.025 545.525 118.755 ;
        RECT  545.825 118.025 546.025 118.755 ;
        RECT  546.32 118.025 546.52 118.755 ;
        RECT  547.14 118.025 547.34 118.755 ;
        RECT  547.635 118.025 547.835 118.755 ;
        RECT  548.135 118.025 548.335 118.755 ;
        RECT  548.29 0.52 548.55 2.335 ;
        RECT  548.635 118.025 548.835 118.755 ;
        RECT  548.8 0.52 549.06 14.11 ;
        RECT  549.13 118.025 549.33 118.755 ;
        RECT  550.175 0.17 550.945 0.94 ;
        RECT  550.685 0.17 550.945 8.7 ;
        RECT  550.175 0.17 550.435 12.9 ;
        RECT  549.665 0.52 549.925 2.485 ;
        RECT  549.95 118.025 550.15 118.755 ;
        RECT  551.195 0.17 551.965 0.43 ;
        RECT  551.705 0.17 551.965 10.48 ;
        RECT  551.195 0.17 551.455 10.99 ;
        RECT  550.445 118.025 550.645 118.755 ;
        RECT  550.945 118.025 551.145 118.755 ;
        RECT  551.445 118.025 551.645 118.755 ;
        RECT  551.94 118.025 552.14 118.755 ;
        RECT  553.235 0.17 554.005 0.43 ;
        RECT  553.235 0.17 553.495 11.5 ;
        RECT  553.745 0.17 554.005 11.5 ;
        RECT  552.76 118.025 552.96 118.755 ;
        RECT  553.255 118.025 553.455 118.755 ;
        RECT  554.255 0.17 555.025 0.94 ;
        RECT  554.255 0.17 554.515 12.9 ;
        RECT  554.765 0.17 555.025 12.9 ;
        RECT  553.755 118.025 553.955 118.755 ;
        RECT  554.255 118.025 554.455 118.755 ;
        RECT  554.75 118.025 554.95 118.755 ;
        RECT  555.275 0.52 555.535 5.815 ;
        RECT  556.13 0.52 556.39 5.16 ;
        RECT  556.13 4.9 556.91 5.16 ;
        RECT  556.65 4.9 556.91 6.64 ;
        RECT  555.57 118.025 555.77 118.755 ;
        RECT  556.065 118.025 556.265 118.755 ;
        RECT  556.565 118.025 556.765 118.755 ;
        RECT  557.065 118.025 557.265 118.755 ;
        RECT  557.56 118.025 557.76 118.755 ;
        RECT  558.38 118.025 558.58 118.755 ;
        RECT  558.875 118.025 559.075 118.755 ;
        RECT  559.375 118.025 559.575 118.755 ;
        RECT  559.53 0.52 559.79 2.335 ;
        RECT  559.875 118.025 560.075 118.755 ;
        RECT  560.04 0.52 560.3 14.11 ;
        RECT  560.37 118.025 560.57 118.755 ;
        RECT  561.415 0.17 562.185 0.94 ;
        RECT  561.925 0.17 562.185 8.7 ;
        RECT  561.415 0.17 561.675 12.9 ;
        RECT  560.905 0.52 561.165 2.485 ;
        RECT  561.19 118.025 561.39 118.755 ;
        RECT  562.435 0.17 563.205 0.43 ;
        RECT  562.945 0.17 563.205 10.48 ;
        RECT  562.435 0.17 562.695 10.99 ;
        RECT  561.685 118.025 561.885 118.755 ;
        RECT  562.185 118.025 562.385 118.755 ;
        RECT  562.685 118.025 562.885 118.755 ;
        RECT  563.18 118.025 563.38 118.755 ;
        RECT  564.475 0.17 565.245 0.43 ;
        RECT  564.475 0.17 564.735 11.5 ;
        RECT  564.985 0.17 565.245 11.5 ;
        RECT  564 118.025 564.2 118.755 ;
        RECT  564.495 118.025 564.695 118.755 ;
        RECT  565.495 0.17 566.265 0.94 ;
        RECT  565.495 0.17 565.755 12.9 ;
        RECT  566.005 0.17 566.265 12.9 ;
        RECT  564.995 118.025 565.195 118.755 ;
        RECT  565.495 118.025 565.695 118.755 ;
        RECT  565.99 118.025 566.19 118.755 ;
        RECT  566.515 0.52 566.775 5.815 ;
        RECT  567.37 0.52 567.63 5.16 ;
        RECT  567.37 4.9 568.15 5.16 ;
        RECT  567.89 4.9 568.15 6.64 ;
        RECT  566.81 118.025 567.01 118.755 ;
        RECT  567.305 118.025 567.505 118.755 ;
        RECT  567.805 118.025 568.005 118.755 ;
        RECT  568.305 118.025 568.505 118.755 ;
        RECT  568.8 118.025 569 118.755 ;
        RECT  569.62 118.025 569.82 118.755 ;
        RECT  570.115 118.025 570.315 118.755 ;
        RECT  570.615 118.025 570.815 118.755 ;
        RECT  570.77 0.52 571.03 2.335 ;
        RECT  571.115 118.025 571.315 118.755 ;
        RECT  571.28 0.52 571.54 14.11 ;
        RECT  571.61 118.025 571.81 118.755 ;
        RECT  572.655 0.17 573.425 0.94 ;
        RECT  573.165 0.17 573.425 8.7 ;
        RECT  572.655 0.17 572.915 12.9 ;
        RECT  572.145 0.52 572.405 2.485 ;
        RECT  572.43 118.025 572.63 118.755 ;
        RECT  573.675 0.17 574.445 0.43 ;
        RECT  574.185 0.17 574.445 10.48 ;
        RECT  573.675 0.17 573.935 10.99 ;
        RECT  572.925 118.025 573.125 118.755 ;
        RECT  573.425 118.025 573.625 118.755 ;
        RECT  573.925 118.025 574.125 118.755 ;
        RECT  574.42 118.025 574.62 118.755 ;
        RECT  575.715 0.17 576.485 0.43 ;
        RECT  575.715 0.17 575.975 11.5 ;
        RECT  576.225 0.17 576.485 11.5 ;
        RECT  575.24 118.025 575.44 118.755 ;
        RECT  575.735 118.025 575.935 118.755 ;
        RECT  576.735 0.17 577.505 0.94 ;
        RECT  576.735 0.17 576.995 12.9 ;
        RECT  577.245 0.17 577.505 12.9 ;
        RECT  576.235 118.025 576.435 118.755 ;
        RECT  576.735 118.025 576.935 118.755 ;
        RECT  577.23 118.025 577.43 118.755 ;
        RECT  577.755 0.52 578.015 5.815 ;
        RECT  578.61 0.52 578.87 5.16 ;
        RECT  578.61 4.9 579.39 5.16 ;
        RECT  579.13 4.9 579.39 6.64 ;
        RECT  578.05 118.025 578.25 118.755 ;
        RECT  578.545 118.025 578.745 118.755 ;
        RECT  579.045 118.025 579.245 118.755 ;
        RECT  579.545 118.025 579.745 118.755 ;
        RECT  580.04 118.025 580.24 118.755 ;
        RECT  580.86 118.025 581.06 118.755 ;
        RECT  581.355 118.025 581.555 118.755 ;
        RECT  581.855 118.025 582.055 118.755 ;
        RECT  582.01 0.52 582.27 2.335 ;
        RECT  582.355 118.025 582.555 118.755 ;
        RECT  582.52 0.52 582.78 14.11 ;
        RECT  582.85 118.025 583.05 118.755 ;
        RECT  583.895 0.17 584.665 0.94 ;
        RECT  584.405 0.17 584.665 8.7 ;
        RECT  583.895 0.17 584.155 12.9 ;
        RECT  583.385 0.52 583.645 2.485 ;
        RECT  583.67 118.025 583.87 118.755 ;
        RECT  584.915 0.17 585.685 0.43 ;
        RECT  585.425 0.17 585.685 10.48 ;
        RECT  584.915 0.17 585.175 10.99 ;
        RECT  584.165 118.025 584.365 118.755 ;
        RECT  584.665 118.025 584.865 118.755 ;
        RECT  585.165 118.025 585.365 118.755 ;
        RECT  585.66 118.025 585.86 118.755 ;
        RECT  586.955 0.17 587.725 0.43 ;
        RECT  586.955 0.17 587.215 11.5 ;
        RECT  587.465 0.17 587.725 11.5 ;
        RECT  586.48 118.025 586.68 118.755 ;
        RECT  586.975 118.025 587.175 118.755 ;
        RECT  587.975 0.17 588.745 0.94 ;
        RECT  587.975 0.17 588.235 12.9 ;
        RECT  588.485 0.17 588.745 12.9 ;
        RECT  587.475 118.025 587.675 118.755 ;
        RECT  587.975 118.025 588.175 118.755 ;
        RECT  588.47 118.025 588.67 118.755 ;
        RECT  588.995 0.52 589.255 5.815 ;
        RECT  589.85 0.52 590.11 5.16 ;
        RECT  589.85 4.9 590.63 5.16 ;
        RECT  590.37 4.9 590.63 6.64 ;
        RECT  589.29 118.025 589.49 118.755 ;
        RECT  589.785 118.025 589.985 118.755 ;
        RECT  590.285 118.025 590.485 118.755 ;
        RECT  590.785 118.025 590.985 118.755 ;
        RECT  591.28 118.025 591.48 118.755 ;
        RECT  592.1 118.025 592.3 118.755 ;
        RECT  592.595 118.025 592.795 118.755 ;
        RECT  593.095 118.025 593.295 118.755 ;
        RECT  593.25 0.52 593.51 2.335 ;
        RECT  593.595 118.025 593.795 118.755 ;
        RECT  593.76 0.52 594.02 14.11 ;
        RECT  594.09 118.025 594.29 118.755 ;
        RECT  595.135 0.17 595.905 0.94 ;
        RECT  595.645 0.17 595.905 8.7 ;
        RECT  595.135 0.17 595.395 12.9 ;
        RECT  594.625 0.52 594.885 2.485 ;
        RECT  594.91 118.025 595.11 118.755 ;
        RECT  596.155 0.17 596.925 0.43 ;
        RECT  596.665 0.17 596.925 10.48 ;
        RECT  596.155 0.17 596.415 10.99 ;
        RECT  595.405 118.025 595.605 118.755 ;
        RECT  595.905 118.025 596.105 118.755 ;
        RECT  596.405 118.025 596.605 118.755 ;
        RECT  596.9 118.025 597.1 118.755 ;
        RECT  598.195 0.17 598.965 0.43 ;
        RECT  598.195 0.17 598.455 11.5 ;
        RECT  598.705 0.17 598.965 11.5 ;
        RECT  597.72 118.025 597.92 118.755 ;
        RECT  598.215 118.025 598.415 118.755 ;
        RECT  599.215 0.17 599.985 0.94 ;
        RECT  599.215 0.17 599.475 12.9 ;
        RECT  599.725 0.17 599.985 12.9 ;
        RECT  598.715 118.025 598.915 118.755 ;
        RECT  599.215 118.025 599.415 118.755 ;
        RECT  599.71 118.025 599.91 118.755 ;
        RECT  600.235 0.52 600.495 5.815 ;
        RECT  601.09 0.52 601.35 5.16 ;
        RECT  601.09 4.9 601.87 5.16 ;
        RECT  601.61 4.9 601.87 6.64 ;
        RECT  600.53 118.025 600.73 118.755 ;
        RECT  601.025 118.025 601.225 118.755 ;
        RECT  601.525 118.025 601.725 118.755 ;
        RECT  602.025 118.025 602.225 118.755 ;
        RECT  602.52 118.025 602.72 118.755 ;
        RECT  603.34 118.025 603.54 118.755 ;
        RECT  603.835 118.025 604.035 118.755 ;
        RECT  604.335 118.025 604.535 118.755 ;
        RECT  604.49 0.52 604.75 2.335 ;
        RECT  604.835 118.025 605.035 118.755 ;
        RECT  605 0.52 605.26 14.11 ;
        RECT  605.33 118.025 605.53 118.755 ;
        RECT  606.375 0.17 607.145 0.94 ;
        RECT  606.885 0.17 607.145 8.7 ;
        RECT  606.375 0.17 606.635 12.9 ;
        RECT  605.865 0.52 606.125 2.485 ;
        RECT  606.15 118.025 606.35 118.755 ;
        RECT  607.395 0.17 608.165 0.43 ;
        RECT  607.905 0.17 608.165 10.48 ;
        RECT  607.395 0.17 607.655 10.99 ;
        RECT  606.645 118.025 606.845 118.755 ;
        RECT  607.145 118.025 607.345 118.755 ;
        RECT  607.645 118.025 607.845 118.755 ;
        RECT  608.14 118.025 608.34 118.755 ;
        RECT  609.435 0.17 610.205 0.43 ;
        RECT  609.435 0.17 609.695 11.5 ;
        RECT  609.945 0.17 610.205 11.5 ;
        RECT  608.96 118.025 609.16 118.755 ;
        RECT  609.455 118.025 609.655 118.755 ;
        RECT  610.455 0.17 611.225 0.94 ;
        RECT  610.455 0.17 610.715 12.9 ;
        RECT  610.965 0.17 611.225 12.9 ;
        RECT  609.955 118.025 610.155 118.755 ;
        RECT  610.455 118.025 610.655 118.755 ;
        RECT  610.95 118.025 611.15 118.755 ;
        RECT  611.475 0.52 611.735 5.815 ;
        RECT  612.33 0.52 612.59 5.16 ;
        RECT  612.33 4.9 613.11 5.16 ;
        RECT  612.85 4.9 613.11 6.64 ;
        RECT  611.77 118.025 611.97 118.755 ;
        RECT  612.265 118.025 612.465 118.755 ;
        RECT  612.765 118.025 612.965 118.755 ;
        RECT  613.265 118.025 613.465 118.755 ;
        RECT  613.76 118.025 613.96 118.755 ;
        RECT  614.58 118.025 614.78 118.755 ;
        RECT  615.075 118.025 615.275 118.755 ;
        RECT  615.575 118.025 615.775 118.755 ;
        RECT  615.73 0.52 615.99 2.335 ;
        RECT  616.075 118.025 616.275 118.755 ;
        RECT  616.24 0.52 616.5 14.11 ;
        RECT  616.57 118.025 616.77 118.755 ;
        RECT  617.615 0.17 618.385 0.94 ;
        RECT  618.125 0.17 618.385 8.7 ;
        RECT  617.615 0.17 617.875 12.9 ;
        RECT  617.105 0.52 617.365 2.485 ;
        RECT  617.39 118.025 617.59 118.755 ;
        RECT  618.635 0.17 619.405 0.43 ;
        RECT  619.145 0.17 619.405 10.48 ;
        RECT  618.635 0.17 618.895 10.99 ;
        RECT  617.885 118.025 618.085 118.755 ;
        RECT  618.385 118.025 618.585 118.755 ;
        RECT  618.885 118.025 619.085 118.755 ;
        RECT  619.38 118.025 619.58 118.755 ;
        RECT  620.675 0.17 621.445 0.43 ;
        RECT  620.675 0.17 620.935 11.5 ;
        RECT  621.185 0.17 621.445 11.5 ;
        RECT  620.2 118.025 620.4 118.755 ;
        RECT  620.695 118.025 620.895 118.755 ;
        RECT  621.695 0.17 622.465 0.94 ;
        RECT  621.695 0.17 621.955 12.9 ;
        RECT  622.205 0.17 622.465 12.9 ;
        RECT  621.195 118.025 621.395 118.755 ;
        RECT  621.695 118.025 621.895 118.755 ;
        RECT  622.19 118.025 622.39 118.755 ;
        RECT  622.715 0.52 622.975 5.815 ;
        RECT  623.57 0.52 623.83 5.16 ;
        RECT  623.57 4.9 624.35 5.16 ;
        RECT  624.09 4.9 624.35 6.64 ;
        RECT  623.01 118.025 623.21 118.755 ;
        RECT  623.505 118.025 623.705 118.755 ;
        RECT  624.005 118.025 624.205 118.755 ;
        RECT  624.505 118.025 624.705 118.755 ;
        RECT  625 118.025 625.2 118.755 ;
        RECT  625.82 118.025 626.02 118.755 ;
        RECT  626.315 118.025 626.515 118.755 ;
        RECT  626.815 118.025 627.015 118.755 ;
        RECT  626.97 0.52 627.23 2.335 ;
        RECT  627.315 118.025 627.515 118.755 ;
        RECT  627.48 0.52 627.74 14.11 ;
        RECT  627.81 118.025 628.01 118.755 ;
        RECT  628.855 0.17 629.625 0.94 ;
        RECT  629.365 0.17 629.625 8.7 ;
        RECT  628.855 0.17 629.115 12.9 ;
        RECT  628.345 0.52 628.605 2.485 ;
        RECT  628.63 118.025 628.83 118.755 ;
        RECT  629.875 0.17 630.645 0.43 ;
        RECT  630.385 0.17 630.645 10.48 ;
        RECT  629.875 0.17 630.135 10.99 ;
        RECT  629.125 118.025 629.325 118.755 ;
        RECT  629.625 118.025 629.825 118.755 ;
        RECT  630.125 118.025 630.325 118.755 ;
        RECT  630.62 118.025 630.82 118.755 ;
        RECT  631.915 0.17 632.685 0.43 ;
        RECT  631.915 0.17 632.175 11.5 ;
        RECT  632.425 0.17 632.685 11.5 ;
        RECT  631.44 118.025 631.64 118.755 ;
        RECT  631.935 118.025 632.135 118.755 ;
        RECT  632.935 0.17 633.705 0.94 ;
        RECT  632.935 0.17 633.195 12.9 ;
        RECT  633.445 0.17 633.705 12.9 ;
        RECT  632.435 118.025 632.635 118.755 ;
        RECT  632.935 118.025 633.135 118.755 ;
        RECT  633.43 118.025 633.63 118.755 ;
        RECT  633.955 0.52 634.215 5.815 ;
        RECT  634.81 0.52 635.07 5.16 ;
        RECT  634.81 4.9 635.59 5.16 ;
        RECT  635.33 4.9 635.59 6.64 ;
        RECT  634.25 118.025 634.45 118.755 ;
        RECT  634.745 118.025 634.945 118.755 ;
        RECT  635.245 118.025 635.445 118.755 ;
        RECT  635.745 118.025 635.945 118.755 ;
        RECT  636.24 118.025 636.44 118.755 ;
        RECT  637.06 118.025 637.26 118.755 ;
        RECT  637.555 118.025 637.755 118.755 ;
        RECT  638.055 118.025 638.255 118.755 ;
        RECT  638.21 0.52 638.47 2.335 ;
        RECT  638.555 118.025 638.755 118.755 ;
        RECT  638.72 0.52 638.98 14.11 ;
        RECT  639.05 118.025 639.25 118.755 ;
        RECT  640.095 0.17 640.865 0.94 ;
        RECT  640.605 0.17 640.865 8.7 ;
        RECT  640.095 0.17 640.355 12.9 ;
        RECT  639.585 0.52 639.845 2.485 ;
        RECT  639.87 118.025 640.07 118.755 ;
        RECT  641.115 0.17 641.885 0.43 ;
        RECT  641.625 0.17 641.885 10.48 ;
        RECT  641.115 0.17 641.375 10.99 ;
        RECT  640.365 118.025 640.565 118.755 ;
        RECT  640.865 118.025 641.065 118.755 ;
        RECT  641.365 118.025 641.565 118.755 ;
        RECT  641.86 118.025 642.06 118.755 ;
        RECT  643.155 0.17 643.925 0.43 ;
        RECT  643.155 0.17 643.415 11.5 ;
        RECT  643.665 0.17 643.925 11.5 ;
        RECT  642.68 118.025 642.88 118.755 ;
        RECT  643.175 118.025 643.375 118.755 ;
        RECT  644.175 0.17 644.945 0.94 ;
        RECT  644.175 0.17 644.435 12.9 ;
        RECT  644.685 0.17 644.945 12.9 ;
        RECT  643.675 118.025 643.875 118.755 ;
        RECT  644.175 118.025 644.375 118.755 ;
        RECT  644.67 118.025 644.87 118.755 ;
        RECT  645.195 0.52 645.455 5.815 ;
        RECT  646.05 0.52 646.31 5.16 ;
        RECT  646.05 4.9 646.83 5.16 ;
        RECT  646.57 4.9 646.83 6.64 ;
        RECT  645.49 118.025 645.69 118.755 ;
        RECT  645.985 118.025 646.185 118.755 ;
        RECT  646.485 118.025 646.685 118.755 ;
        RECT  646.985 118.025 647.185 118.755 ;
        RECT  647.48 118.025 647.68 118.755 ;
        RECT  648.3 118.025 648.5 118.755 ;
        RECT  648.795 118.025 648.995 118.755 ;
        RECT  649.295 118.025 649.495 118.755 ;
        RECT  649.45 0.52 649.71 2.335 ;
        RECT  649.795 118.025 649.995 118.755 ;
        RECT  649.96 0.52 650.22 14.11 ;
        RECT  650.29 118.025 650.49 118.755 ;
        RECT  651.335 0.17 652.105 0.94 ;
        RECT  651.845 0.17 652.105 8.7 ;
        RECT  651.335 0.17 651.595 12.9 ;
        RECT  650.825 0.52 651.085 2.485 ;
        RECT  651.11 118.025 651.31 118.755 ;
        RECT  652.355 0.17 653.125 0.43 ;
        RECT  652.865 0.17 653.125 10.48 ;
        RECT  652.355 0.17 652.615 10.99 ;
        RECT  651.605 118.025 651.805 118.755 ;
        RECT  652.105 118.025 652.305 118.755 ;
        RECT  652.605 118.025 652.805 118.755 ;
        RECT  653.1 118.025 653.3 118.755 ;
        RECT  654.395 0.17 655.165 0.43 ;
        RECT  654.395 0.17 654.655 11.5 ;
        RECT  654.905 0.17 655.165 11.5 ;
        RECT  653.92 118.025 654.12 118.755 ;
        RECT  654.415 118.025 654.615 118.755 ;
        RECT  655.415 0.17 656.185 0.94 ;
        RECT  655.415 0.17 655.675 12.9 ;
        RECT  655.925 0.17 656.185 12.9 ;
        RECT  654.915 118.025 655.115 118.755 ;
        RECT  655.415 118.025 655.615 118.755 ;
        RECT  655.91 118.025 656.11 118.755 ;
        RECT  656.435 0.52 656.695 5.815 ;
        RECT  657.29 0.52 657.55 5.16 ;
        RECT  657.29 4.9 658.07 5.16 ;
        RECT  657.81 4.9 658.07 6.64 ;
        RECT  656.73 118.025 656.93 118.755 ;
        RECT  657.225 118.025 657.425 118.755 ;
        RECT  657.725 118.025 657.925 118.755 ;
        RECT  658.225 118.025 658.425 118.755 ;
        RECT  658.72 118.025 658.92 118.755 ;
        RECT  659.54 118.025 659.74 118.755 ;
        RECT  660.035 118.025 660.235 118.755 ;
        RECT  660.535 118.025 660.735 118.755 ;
        RECT  660.69 0.52 660.95 2.335 ;
        RECT  661.035 118.025 661.235 118.755 ;
        RECT  661.2 0.52 661.46 14.11 ;
        RECT  661.53 118.025 661.73 118.755 ;
        RECT  662.575 0.17 663.345 0.94 ;
        RECT  663.085 0.17 663.345 8.7 ;
        RECT  662.575 0.17 662.835 12.9 ;
        RECT  662.065 0.52 662.325 2.485 ;
        RECT  662.35 118.025 662.55 118.755 ;
        RECT  663.595 0.17 664.365 0.43 ;
        RECT  664.105 0.17 664.365 10.48 ;
        RECT  663.595 0.17 663.855 10.99 ;
        RECT  662.845 118.025 663.045 118.755 ;
        RECT  663.345 118.025 663.545 118.755 ;
        RECT  663.845 118.025 664.045 118.755 ;
        RECT  664.34 118.025 664.54 118.755 ;
        RECT  665.635 0.17 666.405 0.43 ;
        RECT  665.635 0.17 665.895 11.5 ;
        RECT  666.145 0.17 666.405 11.5 ;
        RECT  665.16 118.025 665.36 118.755 ;
        RECT  665.655 118.025 665.855 118.755 ;
        RECT  666.655 0.17 667.425 0.94 ;
        RECT  666.655 0.17 666.915 12.9 ;
        RECT  667.165 0.17 667.425 12.9 ;
        RECT  666.155 118.025 666.355 118.755 ;
        RECT  666.655 118.025 666.855 118.755 ;
        RECT  667.15 118.025 667.35 118.755 ;
        RECT  667.675 0.52 667.935 5.815 ;
        RECT  668.53 0.52 668.79 5.16 ;
        RECT  668.53 4.9 669.31 5.16 ;
        RECT  669.05 4.9 669.31 6.64 ;
        RECT  667.97 118.025 668.17 118.755 ;
        RECT  668.465 118.025 668.665 118.755 ;
        RECT  668.965 118.025 669.165 118.755 ;
        RECT  669.465 118.025 669.665 118.755 ;
        RECT  669.96 118.025 670.16 118.755 ;
        RECT  670.78 118.025 670.98 118.755 ;
        RECT  671.275 118.025 671.475 118.755 ;
        RECT  671.775 118.025 671.975 118.755 ;
        RECT  671.93 0.52 672.19 2.335 ;
        RECT  672.275 118.025 672.475 118.755 ;
        RECT  672.44 0.52 672.7 14.11 ;
        RECT  672.77 118.025 672.97 118.755 ;
        RECT  673.815 0.17 674.585 0.94 ;
        RECT  674.325 0.17 674.585 8.7 ;
        RECT  673.815 0.17 674.075 12.9 ;
        RECT  673.305 0.52 673.565 2.485 ;
        RECT  673.59 118.025 673.79 118.755 ;
        RECT  674.835 0.17 675.605 0.43 ;
        RECT  675.345 0.17 675.605 10.48 ;
        RECT  674.835 0.17 675.095 10.99 ;
        RECT  674.085 118.025 674.285 118.755 ;
        RECT  674.585 118.025 674.785 118.755 ;
        RECT  675.085 118.025 675.285 118.755 ;
        RECT  675.58 118.025 675.78 118.755 ;
        RECT  676.875 0.17 677.645 0.43 ;
        RECT  676.875 0.17 677.135 11.5 ;
        RECT  677.385 0.17 677.645 11.5 ;
        RECT  676.4 118.025 676.6 118.755 ;
        RECT  676.895 118.025 677.095 118.755 ;
        RECT  677.895 0.17 678.665 0.94 ;
        RECT  677.895 0.17 678.155 12.9 ;
        RECT  678.405 0.17 678.665 12.9 ;
        RECT  677.395 118.025 677.595 118.755 ;
        RECT  677.895 118.025 678.095 118.755 ;
        RECT  678.39 118.025 678.59 118.755 ;
        RECT  678.915 0.52 679.175 5.815 ;
        RECT  679.77 0.52 680.03 5.16 ;
        RECT  679.77 4.9 680.55 5.16 ;
        RECT  680.29 4.9 680.55 6.64 ;
        RECT  679.21 118.025 679.41 118.755 ;
        RECT  679.705 118.025 679.905 118.755 ;
        RECT  680.205 118.025 680.405 118.755 ;
        RECT  680.705 118.025 680.905 118.755 ;
        RECT  681.2 118.025 681.4 118.755 ;
        RECT  682.02 118.025 682.22 118.755 ;
        RECT  682.515 118.025 682.715 118.755 ;
        RECT  683.015 118.025 683.215 118.755 ;
        RECT  683.17 0.52 683.43 2.335 ;
        RECT  683.515 118.025 683.715 118.755 ;
        RECT  683.68 0.52 683.94 14.11 ;
        RECT  684.01 118.025 684.21 118.755 ;
        RECT  685.055 0.17 685.825 0.94 ;
        RECT  685.565 0.17 685.825 8.7 ;
        RECT  685.055 0.17 685.315 12.9 ;
        RECT  684.545 0.52 684.805 2.485 ;
        RECT  684.83 118.025 685.03 118.755 ;
        RECT  686.075 0.17 686.845 0.43 ;
        RECT  686.585 0.17 686.845 10.48 ;
        RECT  686.075 0.17 686.335 10.99 ;
        RECT  685.325 118.025 685.525 118.755 ;
        RECT  685.825 118.025 686.025 118.755 ;
        RECT  686.325 118.025 686.525 118.755 ;
        RECT  686.82 118.025 687.02 118.755 ;
        RECT  688.115 0.17 688.885 0.43 ;
        RECT  688.115 0.17 688.375 11.5 ;
        RECT  688.625 0.17 688.885 11.5 ;
        RECT  687.64 118.025 687.84 118.755 ;
        RECT  688.135 118.025 688.335 118.755 ;
        RECT  689.135 0.17 689.905 0.94 ;
        RECT  689.135 0.17 689.395 12.9 ;
        RECT  689.645 0.17 689.905 12.9 ;
        RECT  688.635 118.025 688.835 118.755 ;
        RECT  689.135 118.025 689.335 118.755 ;
        RECT  689.63 118.025 689.83 118.755 ;
        RECT  690.155 0.52 690.415 5.815 ;
        RECT  691.01 0.52 691.27 5.16 ;
        RECT  691.01 4.9 691.79 5.16 ;
        RECT  691.53 4.9 691.79 6.64 ;
        RECT  690.45 118.025 690.65 118.755 ;
        RECT  690.945 118.025 691.145 118.755 ;
        RECT  691.445 118.025 691.645 118.755 ;
        RECT  691.945 118.025 692.145 118.755 ;
        RECT  692.44 118.025 692.64 118.755 ;
        RECT  693.26 118.025 693.46 118.755 ;
        RECT  693.755 118.025 693.955 118.755 ;
        RECT  694.255 118.025 694.455 118.755 ;
        RECT  694.41 0.52 694.67 2.335 ;
        RECT  694.755 118.025 694.955 118.755 ;
        RECT  694.92 0.52 695.18 14.11 ;
        RECT  695.25 118.025 695.45 118.755 ;
        RECT  696.295 0.17 697.065 0.94 ;
        RECT  696.805 0.17 697.065 8.7 ;
        RECT  696.295 0.17 696.555 12.9 ;
        RECT  695.785 0.52 696.045 2.485 ;
        RECT  696.07 118.025 696.27 118.755 ;
        RECT  697.315 0.17 698.085 0.43 ;
        RECT  697.825 0.17 698.085 10.48 ;
        RECT  697.315 0.17 697.575 10.99 ;
        RECT  696.565 118.025 696.765 118.755 ;
        RECT  697.065 118.025 697.265 118.755 ;
        RECT  697.565 118.025 697.765 118.755 ;
        RECT  698.06 118.025 698.26 118.755 ;
        RECT  699.355 0.17 700.125 0.43 ;
        RECT  699.355 0.17 699.615 11.5 ;
        RECT  699.865 0.17 700.125 11.5 ;
        RECT  698.88 118.025 699.08 118.755 ;
        RECT  699.375 118.025 699.575 118.755 ;
        RECT  700.375 0.17 701.145 0.94 ;
        RECT  700.375 0.17 700.635 12.9 ;
        RECT  700.885 0.17 701.145 12.9 ;
        RECT  699.875 118.025 700.075 118.755 ;
        RECT  700.375 118.025 700.575 118.755 ;
        RECT  700.87 118.025 701.07 118.755 ;
        RECT  701.395 0.52 701.655 5.815 ;
        RECT  702.25 0.52 702.51 5.16 ;
        RECT  702.25 4.9 703.03 5.16 ;
        RECT  702.77 4.9 703.03 6.64 ;
        RECT  701.69 118.025 701.89 118.755 ;
        RECT  702.185 118.025 702.385 118.755 ;
        RECT  702.685 118.025 702.885 118.755 ;
        RECT  703.185 118.025 703.385 118.755 ;
        RECT  703.68 118.025 703.88 118.755 ;
        RECT  704.5 118.025 704.7 118.755 ;
        RECT  704.995 118.025 705.195 118.755 ;
        RECT  705.495 118.025 705.695 118.755 ;
        RECT  705.65 0.52 705.91 2.335 ;
        RECT  705.995 118.025 706.195 118.755 ;
        RECT  706.16 0.52 706.42 14.11 ;
        RECT  706.49 118.025 706.69 118.755 ;
        RECT  707.535 0.17 708.305 0.94 ;
        RECT  708.045 0.17 708.305 8.7 ;
        RECT  707.535 0.17 707.795 12.9 ;
        RECT  707.025 0.52 707.285 2.485 ;
        RECT  707.31 118.025 707.51 118.755 ;
        RECT  708.555 0.17 709.325 0.43 ;
        RECT  709.065 0.17 709.325 10.48 ;
        RECT  708.555 0.17 708.815 10.99 ;
        RECT  707.805 118.025 708.005 118.755 ;
        RECT  708.305 118.025 708.505 118.755 ;
        RECT  708.805 118.025 709.005 118.755 ;
        RECT  709.3 118.025 709.5 118.755 ;
        RECT  710.595 0.17 711.365 0.43 ;
        RECT  710.595 0.17 710.855 11.5 ;
        RECT  711.105 0.17 711.365 11.5 ;
        RECT  710.12 118.025 710.32 118.755 ;
        RECT  710.615 118.025 710.815 118.755 ;
        RECT  711.615 0.17 712.385 0.94 ;
        RECT  711.615 0.17 711.875 12.9 ;
        RECT  712.125 0.17 712.385 12.9 ;
        RECT  711.115 118.025 711.315 118.755 ;
        RECT  711.615 118.025 711.815 118.755 ;
        RECT  712.11 118.025 712.31 118.755 ;
        RECT  712.635 0.52 712.895 5.815 ;
        RECT  713.49 0.52 713.75 5.16 ;
        RECT  713.49 4.9 714.27 5.16 ;
        RECT  714.01 4.9 714.27 6.64 ;
        RECT  712.93 118.025 713.13 118.755 ;
        RECT  713.425 118.025 713.625 118.755 ;
        RECT  713.925 118.025 714.125 118.755 ;
        RECT  714.425 118.025 714.625 118.755 ;
        RECT  714.92 118.025 715.12 118.755 ;
        RECT  715.74 118.025 715.94 118.755 ;
        RECT  716.235 118.025 716.435 118.755 ;
        RECT  716.735 118.025 716.935 118.755 ;
        RECT  716.89 0.52 717.15 2.335 ;
        RECT  717.235 118.025 717.435 118.755 ;
        RECT  717.4 0.52 717.66 14.11 ;
        RECT  717.73 118.025 717.93 118.755 ;
        RECT  718.775 0.17 719.545 0.94 ;
        RECT  719.285 0.17 719.545 8.7 ;
        RECT  718.775 0.17 719.035 12.9 ;
        RECT  718.265 0.52 718.525 2.485 ;
        RECT  718.55 118.025 718.75 118.755 ;
        RECT  719.795 0.17 720.565 0.43 ;
        RECT  720.305 0.17 720.565 10.48 ;
        RECT  719.795 0.17 720.055 10.99 ;
        RECT  719.045 118.025 719.245 118.755 ;
        RECT  719.545 118.025 719.745 118.755 ;
        RECT  720.045 118.025 720.245 118.755 ;
        RECT  720.54 118.025 720.74 118.755 ;
        RECT  721.835 0.17 722.605 0.43 ;
        RECT  721.835 0.17 722.095 11.5 ;
        RECT  722.345 0.17 722.605 11.5 ;
        RECT  721.36 118.025 721.56 118.755 ;
        RECT  721.855 118.025 722.055 118.755 ;
        RECT  722.855 0.17 723.625 0.94 ;
        RECT  722.855 0.17 723.115 12.9 ;
        RECT  723.365 0.17 723.625 12.9 ;
        RECT  722.355 118.025 722.555 118.755 ;
        RECT  722.855 118.025 723.055 118.755 ;
        RECT  723.35 118.025 723.55 118.755 ;
        RECT  723.875 0.52 724.135 5.815 ;
        RECT  724.73 0.52 724.99 5.16 ;
        RECT  724.73 4.9 725.51 5.16 ;
        RECT  725.25 4.9 725.51 6.64 ;
        RECT  724.17 118.025 724.37 118.755 ;
        RECT  724.665 118.025 724.865 118.755 ;
        RECT  725.165 118.025 725.365 118.755 ;
        RECT  725.665 118.025 725.865 118.755 ;
        RECT  726.16 118.025 726.36 118.755 ;
        RECT  726.98 118.025 727.18 118.755 ;
        RECT  727.475 118.025 727.675 118.755 ;
        RECT  727.975 118.025 728.175 118.755 ;
        RECT  728.13 0.52 728.39 2.335 ;
        RECT  728.475 118.025 728.675 118.755 ;
        RECT  728.64 0.52 728.9 14.11 ;
        RECT  728.97 118.025 729.17 118.755 ;
        RECT  730.015 0.17 730.785 0.94 ;
        RECT  730.525 0.17 730.785 8.7 ;
        RECT  730.015 0.17 730.275 12.9 ;
        RECT  729.505 0.52 729.765 2.485 ;
        RECT  729.79 118.025 729.99 118.755 ;
        RECT  731.035 0.17 731.805 0.43 ;
        RECT  731.545 0.17 731.805 10.48 ;
        RECT  731.035 0.17 731.295 10.99 ;
        RECT  730.285 118.025 730.485 118.755 ;
        RECT  730.785 118.025 730.985 118.755 ;
        RECT  731.285 118.025 731.485 118.755 ;
        RECT  731.78 118.025 731.98 118.755 ;
        RECT  733.075 0.17 733.845 0.43 ;
        RECT  733.075 0.17 733.335 11.5 ;
        RECT  733.585 0.17 733.845 11.5 ;
        RECT  732.6 118.025 732.8 118.755 ;
        RECT  733.095 118.025 733.295 118.755 ;
        RECT  734.095 0.17 734.865 0.94 ;
        RECT  734.095 0.17 734.355 12.9 ;
        RECT  734.605 0.17 734.865 12.9 ;
        RECT  733.595 118.025 733.795 118.755 ;
        RECT  734.095 118.025 734.295 118.755 ;
        RECT  734.59 118.025 734.79 118.755 ;
        RECT  735.115 0.52 735.375 5.815 ;
        RECT  735.97 0.52 736.23 5.16 ;
        RECT  735.97 4.9 736.75 5.16 ;
        RECT  736.49 4.9 736.75 6.64 ;
        RECT  735.41 118.025 735.61 118.755 ;
        RECT  735.905 118.025 736.105 118.755 ;
        RECT  736.405 118.025 736.605 118.755 ;
        RECT  736.905 118.025 737.105 118.755 ;
        RECT  737.4 118.025 737.6 118.755 ;
        RECT  738.22 118.025 738.42 118.755 ;
        RECT  738.715 118.025 738.915 118.755 ;
        RECT  739.215 118.025 739.415 118.755 ;
        RECT  739.37 0.52 739.63 2.335 ;
        RECT  739.715 118.025 739.915 118.755 ;
        RECT  739.88 0.52 740.14 14.11 ;
        RECT  740.21 118.025 740.41 118.755 ;
        RECT  741.255 0.17 742.025 0.94 ;
        RECT  741.765 0.17 742.025 8.7 ;
        RECT  741.255 0.17 741.515 12.9 ;
        RECT  740.745 0.52 741.005 2.485 ;
        RECT  741.03 118.025 741.23 118.755 ;
        RECT  742.275 0.17 743.045 0.43 ;
        RECT  742.785 0.17 743.045 10.48 ;
        RECT  742.275 0.17 742.535 10.99 ;
        RECT  741.525 118.025 741.725 118.755 ;
        RECT  742.025 118.025 742.225 118.755 ;
        RECT  742.525 118.025 742.725 118.755 ;
        RECT  743.02 118.025 743.22 118.755 ;
        RECT  744.315 0.17 745.085 0.43 ;
        RECT  744.315 0.17 744.575 11.5 ;
        RECT  744.825 0.17 745.085 11.5 ;
        RECT  743.84 118.025 744.04 118.755 ;
        RECT  744.335 118.025 744.535 118.755 ;
        RECT  745.335 0.17 746.105 0.94 ;
        RECT  745.335 0.17 745.595 12.9 ;
        RECT  745.845 0.17 746.105 12.9 ;
        RECT  744.835 118.025 745.035 118.755 ;
        RECT  745.335 118.025 745.535 118.755 ;
        RECT  745.83 118.025 746.03 118.755 ;
        RECT  746.355 0.52 746.615 5.815 ;
        RECT  747.21 0.52 747.47 5.16 ;
        RECT  747.21 4.9 747.99 5.16 ;
        RECT  747.73 4.9 747.99 6.64 ;
        RECT  746.65 118.025 746.85 118.755 ;
        RECT  747.145 118.025 747.345 118.755 ;
        RECT  747.645 118.025 747.845 118.755 ;
        RECT  748.145 118.025 748.345 118.755 ;
        RECT  748.64 118.025 748.84 118.755 ;
        RECT  749.46 118.025 749.66 118.755 ;
        RECT  749.955 118.025 750.155 118.755 ;
        RECT  750.455 118.025 750.655 118.755 ;
        RECT  750.61 0.52 750.87 2.335 ;
        RECT  750.955 118.025 751.155 118.755 ;
        RECT  751.12 0.52 751.38 14.11 ;
        RECT  751.45 118.025 751.65 118.755 ;
        RECT  752.495 0.17 753.265 0.94 ;
        RECT  753.005 0.17 753.265 8.7 ;
        RECT  752.495 0.17 752.755 12.9 ;
        RECT  751.985 0.52 752.245 2.485 ;
        RECT  752.27 118.025 752.47 118.755 ;
        RECT  753.515 0.17 754.285 0.43 ;
        RECT  754.025 0.17 754.285 10.48 ;
        RECT  753.515 0.17 753.775 10.99 ;
        RECT  752.765 118.025 752.965 118.755 ;
        RECT  753.265 118.025 753.465 118.755 ;
        RECT  753.765 118.025 753.965 118.755 ;
        RECT  754.26 118.025 754.46 118.755 ;
        RECT  755.555 0.17 756.325 0.43 ;
        RECT  755.555 0.17 755.815 11.5 ;
        RECT  756.065 0.17 756.325 11.5 ;
        RECT  755.08 118.025 755.28 118.755 ;
        RECT  755.575 118.025 755.775 118.755 ;
        RECT  756.575 0.17 757.345 0.94 ;
        RECT  756.575 0.17 756.835 12.9 ;
        RECT  757.085 0.17 757.345 12.9 ;
        RECT  756.075 118.025 756.275 118.755 ;
        RECT  756.575 118.025 756.775 118.755 ;
        RECT  757.07 118.025 757.27 118.755 ;
        RECT  757.595 0.52 757.855 5.815 ;
        RECT  758.45 0.52 758.71 5.16 ;
        RECT  758.45 4.9 759.23 5.16 ;
        RECT  758.97 4.9 759.23 6.64 ;
        RECT  757.89 118.025 758.09 118.755 ;
        RECT  758.385 118.025 758.585 118.755 ;
        RECT  758.885 118.025 759.085 118.755 ;
        RECT  759.385 118.025 759.585 118.755 ;
        RECT  759.88 118.025 760.08 118.755 ;
        RECT  760.7 118.025 760.9 118.755 ;
        RECT  761.195 118.025 761.395 118.755 ;
        RECT  761.695 118.025 761.895 118.755 ;
        RECT  761.85 0.52 762.11 2.335 ;
        RECT  762.195 118.025 762.395 118.755 ;
        RECT  762.36 0.52 762.62 14.11 ;
        RECT  762.69 118.025 762.89 118.755 ;
        RECT  763.735 0.17 764.505 0.94 ;
        RECT  764.245 0.17 764.505 8.7 ;
        RECT  763.735 0.17 763.995 12.9 ;
        RECT  763.225 0.52 763.485 2.485 ;
        RECT  763.51 118.025 763.71 118.755 ;
        RECT  764.755 0.17 765.525 0.43 ;
        RECT  765.265 0.17 765.525 10.48 ;
        RECT  764.755 0.17 765.015 10.99 ;
        RECT  764.005 118.025 764.205 118.755 ;
        RECT  764.505 118.025 764.705 118.755 ;
        RECT  765.005 118.025 765.205 118.755 ;
        RECT  765.5 118.025 765.7 118.755 ;
        RECT  766.795 0.17 767.565 0.43 ;
        RECT  766.795 0.17 767.055 11.5 ;
        RECT  767.305 0.17 767.565 11.5 ;
        RECT  766.32 118.025 766.52 118.755 ;
        RECT  766.815 118.025 767.015 118.755 ;
        RECT  767.815 0.17 768.585 0.94 ;
        RECT  767.815 0.17 768.075 12.9 ;
        RECT  768.325 0.17 768.585 12.9 ;
        RECT  767.315 118.025 767.515 118.755 ;
        RECT  767.815 118.025 768.015 118.755 ;
        RECT  768.31 118.025 768.51 118.755 ;
        RECT  768.835 0.52 769.095 5.815 ;
        RECT  769.69 0.52 769.95 5.16 ;
        RECT  769.69 4.9 770.47 5.16 ;
        RECT  770.21 4.9 770.47 6.64 ;
        RECT  769.13 118.025 769.33 118.755 ;
        RECT  769.625 118.025 769.825 118.755 ;
        RECT  770.125 118.025 770.325 118.755 ;
        RECT  770.625 118.025 770.825 118.755 ;
        RECT  771.12 118.025 771.32 118.755 ;
        RECT  771.94 118.025 772.14 118.755 ;
        RECT  772.435 118.025 772.635 118.755 ;
        RECT  772.935 118.025 773.135 118.755 ;
        RECT  773.09 0.52 773.35 2.335 ;
        RECT  773.435 118.025 773.635 118.755 ;
        RECT  773.6 0.52 773.86 14.11 ;
        RECT  773.93 118.025 774.13 118.755 ;
        RECT  774.975 0.17 775.745 0.94 ;
        RECT  775.485 0.17 775.745 8.7 ;
        RECT  774.975 0.17 775.235 12.9 ;
        RECT  774.465 0.52 774.725 2.485 ;
        RECT  774.75 118.025 774.95 118.755 ;
        RECT  775.995 0.17 776.765 0.43 ;
        RECT  776.505 0.17 776.765 10.48 ;
        RECT  775.995 0.17 776.255 10.99 ;
        RECT  775.245 118.025 775.445 118.755 ;
        RECT  775.745 118.025 775.945 118.755 ;
        RECT  776.245 118.025 776.445 118.755 ;
        RECT  776.74 118.025 776.94 118.755 ;
        RECT  778.035 0.17 778.805 0.43 ;
        RECT  778.035 0.17 778.295 11.5 ;
        RECT  778.545 0.17 778.805 11.5 ;
        RECT  777.56 118.025 777.76 118.755 ;
        RECT  778.055 118.025 778.255 118.755 ;
        RECT  779.055 0.17 779.825 0.94 ;
        RECT  779.055 0.17 779.315 12.9 ;
        RECT  779.565 0.17 779.825 12.9 ;
        RECT  778.555 118.025 778.755 118.755 ;
        RECT  779.055 118.025 779.255 118.755 ;
        RECT  779.55 118.025 779.75 118.755 ;
        RECT  780.075 0.52 780.335 5.815 ;
        RECT  780.93 0.52 781.19 5.16 ;
        RECT  780.93 4.9 781.71 5.16 ;
        RECT  781.45 4.9 781.71 6.64 ;
        RECT  780.37 118.025 780.57 118.755 ;
        RECT  780.865 118.025 781.065 118.755 ;
        RECT  781.365 118.025 781.565 118.755 ;
        RECT  781.865 118.025 782.065 118.755 ;
        RECT  782.36 118.025 782.56 118.755 ;
        RECT  783.18 118.025 783.38 118.755 ;
        RECT  784.175 45.465 784.375 118.755 ;
        RECT  184.505 0 189.335 118.78 ;
        RECT  195.745 0 200.575 118.78 ;
        RECT  206.985 0 211.815 118.78 ;
        RECT  218.225 0 223.055 118.78 ;
        RECT  229.465 0 234.295 118.78 ;
        RECT  240.705 0 245.535 118.78 ;
        RECT  251.945 0 256.775 118.78 ;
        RECT  263.185 0 268.015 118.78 ;
        RECT  274.425 0 279.255 118.78 ;
        RECT  285.665 0 290.495 118.78 ;
        RECT  296.905 0 301.735 118.78 ;
        RECT  308.145 0 312.975 118.78 ;
        RECT  319.385 0 324.215 118.78 ;
        RECT  330.625 0 335.455 118.78 ;
        RECT  341.865 0 346.695 118.78 ;
        RECT  353.105 0 357.935 118.78 ;
        RECT  378.24 0 384.61 118.78 ;
        RECT  393.55 0 394.81 118.78 ;
        RECT  426.545 0 431.375 118.78 ;
        RECT  437.785 0 442.615 118.78 ;
        RECT  449.025 0 453.855 118.78 ;
        RECT  460.265 0 465.095 118.78 ;
        RECT  471.505 0 476.335 118.78 ;
        RECT  482.745 0 487.575 118.78 ;
        RECT  493.985 0 498.815 118.78 ;
        RECT  505.225 0 510.055 118.78 ;
        RECT  516.465 0 521.295 118.78 ;
        RECT  527.705 0 532.535 118.78 ;
        RECT  538.945 0 543.775 118.78 ;
        RECT  550.185 0 555.015 118.78 ;
        RECT  561.425 0 566.255 118.78 ;
        RECT  572.665 0 577.495 118.78 ;
        RECT  583.905 0 588.735 118.78 ;
        RECT  595.145 0 599.975 118.78 ;
        RECT  606.385 0 611.215 118.78 ;
        RECT  617.625 0 622.455 118.78 ;
        RECT  628.865 0 633.695 118.78 ;
        RECT  640.105 0 644.935 118.78 ;
        RECT  651.345 0 656.175 118.78 ;
        RECT  662.585 0 667.415 118.78 ;
        RECT  673.825 0 678.655 118.78 ;
        RECT  685.065 0 689.895 118.78 ;
        RECT  696.305 0 701.135 118.78 ;
        RECT  707.545 0 712.375 118.78 ;
        RECT  718.785 0 723.615 118.78 ;
        RECT  730.025 0 734.855 118.78 ;
        RECT  741.265 0 746.095 118.78 ;
        RECT  752.505 0 757.335 118.78 ;
        RECT  763.745 0 768.575 118.78 ;
        RECT  774.985 0 779.815 118.78 ;
        RECT  385.9 0 386.14 118.78 ;
        RECT  387.43 0 387.67 118.78 ;
        RECT  390.49 0 390.73 118.78 ;
        RECT  392.02 0 392.26 118.78 ;
        RECT  399.15 0 408.07 118.78 ;
        RECT  0 0 3.03 118.78 ;
        RECT  4.655 0.17 9.505 118.78 ;
        RECT  11.65 0 14.27 118.78 ;
        RECT  15.895 0.17 20.745 118.78 ;
        RECT  22.89 0 25.51 118.78 ;
        RECT  27.135 0.17 31.985 118.78 ;
        RECT  34.13 0 36.75 118.78 ;
        RECT  38.375 0.17 43.225 118.78 ;
        RECT  45.37 0 47.99 118.78 ;
        RECT  49.615 0.17 54.465 118.78 ;
        RECT  56.61 0 59.23 118.78 ;
        RECT  60.855 0.17 65.705 118.78 ;
        RECT  67.85 0 70.47 118.78 ;
        RECT  72.095 0.17 76.945 118.78 ;
        RECT  79.09 0 81.71 118.78 ;
        RECT  83.335 0.17 88.185 118.78 ;
        RECT  90.33 0 92.95 118.78 ;
        RECT  94.575 0.17 99.425 118.78 ;
        RECT  101.57 0 104.19 118.78 ;
        RECT  105.815 0.17 110.665 118.78 ;
        RECT  112.81 0 115.43 118.78 ;
        RECT  117.055 0.17 121.905 118.78 ;
        RECT  124.05 0 126.67 118.78 ;
        RECT  128.295 0.17 133.145 118.78 ;
        RECT  135.29 0 137.91 118.78 ;
        RECT  139.535 0.17 144.385 118.78 ;
        RECT  146.53 0 149.15 118.78 ;
        RECT  150.775 0.17 155.625 118.78 ;
        RECT  157.77 0 160.39 118.78 ;
        RECT  162.015 0.17 166.865 118.78 ;
        RECT  169.01 0 171.63 118.78 ;
        RECT  173.255 0.17 178.105 118.78 ;
        RECT  180.25 0 182.87 118.78 ;
        RECT  184.495 0.17 189.345 118.78 ;
        RECT  191.49 0 194.11 118.78 ;
        RECT  195.735 0.17 200.585 118.78 ;
        RECT  202.73 0 205.35 118.78 ;
        RECT  206.975 0.17 211.825 118.78 ;
        RECT  213.97 0 216.59 118.78 ;
        RECT  218.215 0.17 223.065 118.78 ;
        RECT  225.21 0 227.83 118.78 ;
        RECT  229.455 0.17 234.305 118.78 ;
        RECT  236.45 0 239.07 118.78 ;
        RECT  240.695 0.17 245.545 118.78 ;
        RECT  247.69 0 250.31 118.78 ;
        RECT  251.935 0.17 256.785 118.78 ;
        RECT  258.93 0 261.55 118.78 ;
        RECT  263.175 0.17 268.025 118.78 ;
        RECT  270.17 0 272.79 118.78 ;
        RECT  274.415 0.17 279.265 118.78 ;
        RECT  281.41 0 284.03 118.78 ;
        RECT  285.655 0.17 290.505 118.78 ;
        RECT  292.65 0 295.27 118.78 ;
        RECT  296.895 0.17 301.745 118.78 ;
        RECT  303.89 0 306.51 118.78 ;
        RECT  308.135 0.17 312.985 118.78 ;
        RECT  315.13 0 317.75 118.78 ;
        RECT  319.375 0.17 324.225 118.78 ;
        RECT  326.37 0 328.99 118.78 ;
        RECT  330.615 0.17 335.465 118.78 ;
        RECT  337.61 0 340.23 118.78 ;
        RECT  341.855 0.17 346.705 118.78 ;
        RECT  348.85 0 351.47 118.78 ;
        RECT  353.095 0.17 357.945 118.78 ;
        RECT  360.09 0 375.95 118.78 ;
        RECT  378.24 0.17 384.62 118.78 ;
        RECT  385.89 0.3 386.15 118.78 ;
        RECT  387.42 0.3 387.68 118.78 ;
        RECT  390.48 0.3 390.74 118.78 ;
        RECT  392.01 0.3 392.27 118.78 ;
        RECT  393.55 0.17 394.82 118.78 ;
        RECT  393.54 0.3 394.82 118.78 ;
        RECT  399.15 0.3 408.08 118.78 ;
        RECT  408.85 0 424.39 118.78 ;
        RECT  408.84 0.17 424.39 118.78 ;
        RECT  426.535 0.17 431.385 118.78 ;
        RECT  433.01 0 435.63 118.78 ;
        RECT  437.775 0.17 442.625 118.78 ;
        RECT  444.25 0 446.87 118.78 ;
        RECT  449.015 0.17 453.865 118.78 ;
        RECT  455.49 0 458.11 118.78 ;
        RECT  460.255 0.17 465.105 118.78 ;
        RECT  466.73 0 469.35 118.78 ;
        RECT  471.495 0.17 476.345 118.78 ;
        RECT  477.97 0 480.59 118.78 ;
        RECT  482.735 0.17 487.585 118.78 ;
        RECT  489.21 0 491.83 118.78 ;
        RECT  493.975 0.17 498.825 118.78 ;
        RECT  500.45 0 503.07 118.78 ;
        RECT  505.215 0.17 510.065 118.78 ;
        RECT  511.69 0 514.31 118.78 ;
        RECT  516.455 0.17 521.305 118.78 ;
        RECT  522.93 0 525.55 118.78 ;
        RECT  527.695 0.17 532.545 118.78 ;
        RECT  534.17 0 536.79 118.78 ;
        RECT  538.935 0.17 543.785 118.78 ;
        RECT  545.41 0 548.03 118.78 ;
        RECT  550.175 0.17 555.025 118.78 ;
        RECT  556.65 0 559.27 118.78 ;
        RECT  561.415 0.17 566.265 118.78 ;
        RECT  567.89 0 570.51 118.78 ;
        RECT  572.655 0.17 577.505 118.78 ;
        RECT  579.13 0 581.75 118.78 ;
        RECT  583.895 0.17 588.745 118.78 ;
        RECT  590.37 0 592.99 118.78 ;
        RECT  595.135 0.17 599.985 118.78 ;
        RECT  601.61 0 604.23 118.78 ;
        RECT  606.375 0.17 611.225 118.78 ;
        RECT  612.85 0 615.47 118.78 ;
        RECT  617.615 0.17 622.465 118.78 ;
        RECT  624.09 0 626.71 118.78 ;
        RECT  628.855 0.17 633.705 118.78 ;
        RECT  635.33 0 637.95 118.78 ;
        RECT  640.095 0.17 644.945 118.78 ;
        RECT  646.57 0 649.19 118.78 ;
        RECT  651.335 0.17 656.185 118.78 ;
        RECT  657.81 0 660.43 118.78 ;
        RECT  662.575 0.17 667.425 118.78 ;
        RECT  669.05 0 671.67 118.78 ;
        RECT  673.815 0.17 678.665 118.78 ;
        RECT  680.29 0 682.91 118.78 ;
        RECT  685.055 0.17 689.905 118.78 ;
        RECT  691.53 0 694.15 118.78 ;
        RECT  696.295 0.17 701.145 118.78 ;
        RECT  702.77 0 705.39 118.78 ;
        RECT  707.535 0.17 712.385 118.78 ;
        RECT  714.01 0 716.63 118.78 ;
        RECT  718.775 0.17 723.625 118.78 ;
        RECT  725.25 0 727.87 118.78 ;
        RECT  730.015 0.17 734.865 118.78 ;
        RECT  736.49 0 739.11 118.78 ;
        RECT  741.255 0.17 746.105 118.78 ;
        RECT  747.73 0 750.35 118.78 ;
        RECT  752.495 0.17 757.345 118.78 ;
        RECT  758.97 0 761.59 118.78 ;
        RECT  763.735 0.17 768.585 118.78 ;
        RECT  770.21 0 772.83 118.78 ;
        RECT  774.975 0.17 779.825 118.78 ;
        RECT  781.45 0 784.48 118.78 ;
        RECT  0 0.52 784.48 118.78 ;
        RECT  4.665 0 9.495 118.78 ;
        RECT  15.905 0 20.735 118.78 ;
        RECT  27.145 0 31.975 118.78 ;
        RECT  38.385 0 43.215 118.78 ;
        RECT  49.625 0 54.455 118.78 ;
        RECT  60.865 0 65.695 118.78 ;
        RECT  72.105 0 76.935 118.78 ;
        RECT  83.345 0 88.175 118.78 ;
        RECT  94.585 0 99.415 118.78 ;
        RECT  105.825 0 110.655 118.78 ;
        RECT  117.065 0 121.895 118.78 ;
        RECT  128.305 0 133.135 118.78 ;
        RECT  139.545 0 144.375 118.78 ;
        RECT  150.785 0 155.615 118.78 ;
        RECT  162.025 0 166.855 118.78 ;
        RECT  173.265 0 178.095 118.78 ;
      LAYER Metal3 ;
        RECT  0 0 784.48 118.78 ;
      LAYER Metal4 ;
        RECT  0 39.085 9.62 45.205 ;
        RECT  0 0 4 118.78 ;
        RECT  7.33 0 9.62 118.78 ;
        RECT  12.95 39.085 20.86 45.205 ;
        RECT  12.95 0 15.24 118.78 ;
        RECT  18.57 0 20.86 118.78 ;
        RECT  24.19 39.085 32.1 45.205 ;
        RECT  24.19 0 26.48 118.78 ;
        RECT  29.81 0 32.1 118.78 ;
        RECT  35.43 39.085 43.34 45.205 ;
        RECT  35.43 0 37.72 118.78 ;
        RECT  41.05 0 43.34 118.78 ;
        RECT  46.67 39.085 54.58 45.205 ;
        RECT  46.67 0 48.96 118.78 ;
        RECT  52.29 0 54.58 118.78 ;
        RECT  57.91 39.085 65.82 45.205 ;
        RECT  57.91 0 60.2 118.78 ;
        RECT  63.53 0 65.82 118.78 ;
        RECT  69.15 39.085 77.06 45.205 ;
        RECT  69.15 0 71.44 118.78 ;
        RECT  74.77 0 77.06 118.78 ;
        RECT  80.39 39.085 88.3 45.205 ;
        RECT  80.39 0 82.68 118.78 ;
        RECT  86.01 0 88.3 118.78 ;
        RECT  91.63 39.085 99.54 45.205 ;
        RECT  91.63 0 93.92 118.78 ;
        RECT  97.25 0 99.54 118.78 ;
        RECT  102.87 39.085 110.78 45.205 ;
        RECT  102.87 0 105.16 118.78 ;
        RECT  108.49 0 110.78 118.78 ;
        RECT  114.11 39.085 122.02 45.205 ;
        RECT  114.11 0 116.4 118.78 ;
        RECT  119.73 0 122.02 118.78 ;
        RECT  125.35 39.085 133.26 45.205 ;
        RECT  125.35 0 127.64 118.78 ;
        RECT  130.97 0 133.26 118.78 ;
        RECT  136.59 39.085 144.5 45.205 ;
        RECT  136.59 0 138.88 118.78 ;
        RECT  142.21 0 144.5 118.78 ;
        RECT  147.83 39.085 155.74 45.205 ;
        RECT  147.83 0 150.12 118.78 ;
        RECT  153.45 0 155.74 118.78 ;
        RECT  159.07 39.085 166.98 45.205 ;
        RECT  159.07 0 161.36 118.78 ;
        RECT  164.69 0 166.98 118.78 ;
        RECT  170.31 39.085 178.22 45.205 ;
        RECT  170.31 0 172.6 118.78 ;
        RECT  175.93 0 178.22 118.78 ;
        RECT  181.55 39.085 189.46 45.205 ;
        RECT  181.55 0 183.84 118.78 ;
        RECT  187.17 0 189.46 118.78 ;
        RECT  192.79 39.085 200.7 45.205 ;
        RECT  192.79 0 195.08 118.78 ;
        RECT  198.41 0 200.7 118.78 ;
        RECT  204.03 39.085 211.94 45.205 ;
        RECT  204.03 0 206.32 118.78 ;
        RECT  209.65 0 211.94 118.78 ;
        RECT  215.27 39.085 223.18 45.205 ;
        RECT  215.27 0 217.56 118.78 ;
        RECT  220.89 0 223.18 118.78 ;
        RECT  226.51 39.085 234.42 45.205 ;
        RECT  226.51 0 228.8 118.78 ;
        RECT  232.13 0 234.42 118.78 ;
        RECT  237.75 39.085 245.66 45.205 ;
        RECT  237.75 0 240.04 118.78 ;
        RECT  243.37 0 245.66 118.78 ;
        RECT  248.99 39.085 256.9 45.205 ;
        RECT  248.99 0 251.28 118.78 ;
        RECT  254.61 0 256.9 118.78 ;
        RECT  260.23 39.085 268.14 45.205 ;
        RECT  260.23 0 262.52 118.78 ;
        RECT  265.85 0 268.14 118.78 ;
        RECT  271.47 39.085 279.38 45.205 ;
        RECT  271.47 0 273.76 118.78 ;
        RECT  277.09 0 279.38 118.78 ;
        RECT  282.71 39.085 290.62 45.205 ;
        RECT  282.71 0 285 118.78 ;
        RECT  288.33 0 290.62 118.78 ;
        RECT  293.95 39.085 301.86 45.205 ;
        RECT  293.95 0 296.24 118.78 ;
        RECT  299.57 0 301.86 118.78 ;
        RECT  305.19 39.085 313.1 45.205 ;
        RECT  305.19 0 307.48 118.78 ;
        RECT  310.81 0 313.1 118.78 ;
        RECT  316.43 39.085 324.34 45.205 ;
        RECT  316.43 0 318.72 118.78 ;
        RECT  322.05 0 324.34 118.78 ;
        RECT  327.67 39.085 335.58 45.205 ;
        RECT  327.67 0 329.96 118.78 ;
        RECT  333.29 0 335.58 118.78 ;
        RECT  338.91 39.085 346.82 45.205 ;
        RECT  338.91 0 341.2 118.78 ;
        RECT  344.53 0 346.82 118.78 ;
        RECT  350.15 39.085 358.06 45.205 ;
        RECT  350.15 0 352.44 118.78 ;
        RECT  355.77 0 358.06 118.78 ;
        RECT  361.39 0 372.55 118.78 ;
        RECT  375.88 0 377.7 118.78 ;
        RECT  381.03 0 382.85 118.78 ;
        RECT  386.18 0 388 118.78 ;
        RECT  391.33 0 393.15 118.78 ;
        RECT  396.48 0 398.3 118.78 ;
        RECT  426.42 39.085 434.33 45.205 ;
        RECT  426.42 0 428.71 118.78 ;
        RECT  432.04 0 434.33 118.78 ;
        RECT  437.66 39.085 445.57 45.205 ;
        RECT  437.66 0 439.95 118.78 ;
        RECT  443.28 0 445.57 118.78 ;
        RECT  448.9 39.085 456.81 45.205 ;
        RECT  448.9 0 451.19 118.78 ;
        RECT  454.52 0 456.81 118.78 ;
        RECT  460.14 39.085 468.05 45.205 ;
        RECT  460.14 0 462.43 118.78 ;
        RECT  465.76 0 468.05 118.78 ;
        RECT  471.38 39.085 479.29 45.205 ;
        RECT  471.38 0 473.67 118.78 ;
        RECT  477 0 479.29 118.78 ;
        RECT  482.62 39.085 490.53 45.205 ;
        RECT  482.62 0 484.91 118.78 ;
        RECT  488.24 0 490.53 118.78 ;
        RECT  493.86 39.085 501.77 45.205 ;
        RECT  493.86 0 496.15 118.78 ;
        RECT  499.48 0 501.77 118.78 ;
        RECT  505.1 39.085 513.01 45.205 ;
        RECT  505.1 0 507.39 118.78 ;
        RECT  510.72 0 513.01 118.78 ;
        RECT  516.34 39.085 524.25 45.205 ;
        RECT  516.34 0 518.63 118.78 ;
        RECT  521.96 0 524.25 118.78 ;
        RECT  527.58 39.085 535.49 45.205 ;
        RECT  527.58 0 529.87 118.78 ;
        RECT  533.2 0 535.49 118.78 ;
        RECT  538.82 39.085 546.73 45.205 ;
        RECT  538.82 0 541.11 118.78 ;
        RECT  544.44 0 546.73 118.78 ;
        RECT  550.06 39.085 557.97 45.205 ;
        RECT  550.06 0 552.35 118.78 ;
        RECT  555.68 0 557.97 118.78 ;
        RECT  561.3 39.085 569.21 45.205 ;
        RECT  561.3 0 563.59 118.78 ;
        RECT  566.92 0 569.21 118.78 ;
        RECT  572.54 39.085 580.45 45.205 ;
        RECT  572.54 0 574.83 118.78 ;
        RECT  578.16 0 580.45 118.78 ;
        RECT  583.78 39.085 591.69 45.205 ;
        RECT  583.78 0 586.07 118.78 ;
        RECT  589.4 0 591.69 118.78 ;
        RECT  595.02 39.085 602.93 45.205 ;
        RECT  595.02 0 597.31 118.78 ;
        RECT  600.64 0 602.93 118.78 ;
        RECT  606.26 39.085 614.17 45.205 ;
        RECT  606.26 0 608.55 118.78 ;
        RECT  611.88 0 614.17 118.78 ;
        RECT  617.5 39.085 625.41 45.205 ;
        RECT  617.5 0 619.79 118.78 ;
        RECT  623.12 0 625.41 118.78 ;
        RECT  628.74 39.085 636.65 45.205 ;
        RECT  628.74 0 631.03 118.78 ;
        RECT  634.36 0 636.65 118.78 ;
        RECT  639.98 39.085 647.89 45.205 ;
        RECT  639.98 0 642.27 118.78 ;
        RECT  645.6 0 647.89 118.78 ;
        RECT  651.22 39.085 659.13 45.205 ;
        RECT  651.22 0 653.51 118.78 ;
        RECT  656.84 0 659.13 118.78 ;
        RECT  662.46 39.085 670.37 45.205 ;
        RECT  662.46 0 664.75 118.78 ;
        RECT  668.08 0 670.37 118.78 ;
        RECT  673.7 39.085 681.61 45.205 ;
        RECT  673.7 0 675.99 118.78 ;
        RECT  679.32 0 681.61 118.78 ;
        RECT  684.94 39.085 692.85 45.205 ;
        RECT  684.94 0 687.23 118.78 ;
        RECT  690.56 0 692.85 118.78 ;
        RECT  696.18 39.085 704.09 45.205 ;
        RECT  696.18 0 698.47 118.78 ;
        RECT  701.8 0 704.09 118.78 ;
        RECT  707.42 39.085 715.33 45.205 ;
        RECT  707.42 0 709.71 118.78 ;
        RECT  713.04 0 715.33 118.78 ;
        RECT  718.66 39.085 726.57 45.205 ;
        RECT  718.66 0 720.95 118.78 ;
        RECT  724.28 0 726.57 118.78 ;
        RECT  729.9 39.085 737.81 45.205 ;
        RECT  729.9 0 732.19 118.78 ;
        RECT  735.52 0 737.81 118.78 ;
        RECT  741.14 39.085 749.05 45.205 ;
        RECT  741.14 0 743.43 118.78 ;
        RECT  746.76 0 749.05 118.78 ;
        RECT  752.38 39.085 760.29 45.205 ;
        RECT  752.38 0 754.67 118.78 ;
        RECT  758 0 760.29 118.78 ;
        RECT  763.62 39.085 771.53 45.205 ;
        RECT  763.62 0 765.91 118.78 ;
        RECT  769.24 0 771.53 118.78 ;
        RECT  774.86 39.085 784.48 45.205 ;
        RECT  774.86 0 777.15 118.78 ;
        RECT  780.48 0 784.48 118.78 ;
        RECT  401.63 0 403.45 118.78 ;
        RECT  406.78 0 408.6 118.78 ;
        RECT  411.93 0 423.09 118.78 ;
    END
END RM_IHPSG13_1P_256x64_c2_bm_bist
END LIBRARY
