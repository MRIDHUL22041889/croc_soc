VERSION 5.7 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

PROPERTYDEFINITIONS
END PROPERTYDEFINITIONS


MACRO RM_IHPSG13_1P_512x32_c2_bm_bist
    CLASS BLOCK ;
    SIZE 416.64 BY 191.34 ;
    SYMMETRY X Y R90 ;
    PIN A_DIN[16]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  244.49 0 244.75 0.26 ;
        END
    END A_DIN[16]
    PIN A_DIN[15]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  171.89 0 172.15 0.26 ;
        END
    END A_DIN[15]
    PIN A_BIST_DIN[16]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  243.635 0 243.895 0.26 ;
        END
    END A_BIST_DIN[16]
    PIN A_BIST_DIN[15]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  172.745 0 173.005 0.26 ;
        END
    END A_BIST_DIN[15]
    PIN A_BM[16]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  236.65 0 236.91 0.26 ;
        END
    END A_BM[16]
    PIN A_BM[15]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  179.73 0 179.99 0.26 ;
        END
    END A_BM[15]
    PIN A_BIST_BM[16]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  238.025 0 238.285 0.26 ;
        END
    END A_BIST_BM[16]
    PIN A_BIST_BM[15]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  178.355 0 178.615 0.26 ;
        END
    END A_BIST_BM[15]
    PIN A_DOUT[16]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  237.16 0 237.42 0.26 ;
        END
    END A_DOUT[16]
    PIN A_DOUT[15]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  179.22 0 179.48 0.26 ;
        END
    END A_DOUT[15]
    PIN VSS!
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal4 ;
              RECT  403.95 0 406.76 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  392.71 0 395.52 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  381.47 0 384.28 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  370.23 0 373.04 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  358.99 0 361.8 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  347.75 0 350.56 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  336.51 0 339.32 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  325.27 0 328.08 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  314.03 0 316.84 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  302.79 0 305.6 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  291.55 0 294.36 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  280.31 0 283.12 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  269.07 0 271.88 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  257.83 0 260.64 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  246.59 0 249.4 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  235.35 0 238.16 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  224.94 0 227.75 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  214.64 0 217.45 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  199.19 0 202 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  188.89 0 191.7 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  178.48 0 181.29 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  167.24 0 170.05 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  156 0 158.81 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  144.76 0 147.57 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  133.52 0 136.33 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  122.28 0 125.09 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  111.04 0 113.85 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  99.8 0 102.61 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  88.56 0 91.37 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  77.32 0 80.13 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  66.08 0 68.89 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  54.84 0 57.65 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  43.6 0 46.41 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  32.36 0 35.17 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  21.12 0 23.93 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  9.88 0 12.69 191.34 ;
        END
    END VSS!
    PIN VDD!
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal4 ;
              RECT  409.57 0 412.38 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  398.33 0 401.14 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  387.09 0 389.9 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  375.85 0 378.66 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  364.61 0 367.42 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  353.37 0 356.18 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  342.13 0 344.94 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  330.89 0 333.7 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  319.65 0 322.46 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  308.41 0 311.22 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  297.17 0 299.98 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  285.93 0 288.74 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  274.69 0 277.5 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  263.45 0 266.26 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  252.21 0 255.02 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  240.97 0 243.78 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  219.79 0 222.6 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  209.49 0 212.3 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  204.34 0 207.15 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  194.04 0 196.85 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  172.86 0 175.67 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  161.62 0 164.43 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  150.38 0 153.19 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  139.14 0 141.95 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  127.9 0 130.71 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  116.66 0 119.47 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  105.42 0 108.23 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  94.18 0 96.99 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  82.94 0 85.75 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  71.7 0 74.51 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  60.46 0 63.27 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  49.22 0 52.03 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  37.98 0 40.79 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  26.74 0 29.55 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  15.5 0 18.31 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  4.26 0 7.07 38.825 ;
        END
    END VDD!
    PIN VDDARRAY!
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal4 ;
              RECT  409.57 45.465 412.38 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  398.33 45.465 401.14 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  387.09 45.465 389.9 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  375.85 45.465 378.66 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  364.61 45.465 367.42 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  353.37 45.465 356.18 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  342.13 45.465 344.94 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  330.89 45.465 333.7 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  319.65 45.465 322.46 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  308.41 45.465 311.22 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  297.17 45.465 299.98 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  285.93 45.465 288.74 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  274.69 45.465 277.5 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  263.45 45.465 266.26 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  252.21 45.465 255.02 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  240.97 45.465 243.78 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  172.86 45.465 175.67 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  161.62 45.465 164.43 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  150.38 45.465 153.19 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  139.14 45.465 141.95 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  127.9 45.465 130.71 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  116.66 45.465 119.47 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  105.42 45.465 108.23 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  94.18 45.465 96.99 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  82.94 45.465 85.75 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  71.7 45.465 74.51 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  60.46 45.465 63.27 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  49.22 45.465 52.03 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  37.98 45.465 40.79 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  26.74 45.465 29.55 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  15.5 45.465 18.31 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  4.26 45.465 7.07 191.34 ;
        END
    END VDDARRAY!
    PIN A_DIN[17]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  255.73 0 255.99 0.26 ;
        END
    END A_DIN[17]
    PIN A_DIN[14]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  160.65 0 160.91 0.26 ;
        END
    END A_DIN[14]
    PIN A_BIST_DIN[17]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  254.875 0 255.135 0.26 ;
        END
    END A_BIST_DIN[17]
    PIN A_BIST_DIN[14]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  161.505 0 161.765 0.26 ;
        END
    END A_BIST_DIN[14]
    PIN A_BM[17]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  247.89 0 248.15 0.26 ;
        END
    END A_BM[17]
    PIN A_BM[14]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  168.49 0 168.75 0.26 ;
        END
    END A_BM[14]
    PIN A_BIST_BM[17]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  249.265 0 249.525 0.26 ;
        END
    END A_BIST_BM[17]
    PIN A_BIST_BM[14]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  167.115 0 167.375 0.26 ;
        END
    END A_BIST_BM[14]
    PIN A_DOUT[17]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  248.4 0 248.66 0.26 ;
        END
    END A_DOUT[17]
    PIN A_DOUT[14]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  167.98 0 168.24 0.26 ;
        END
    END A_DOUT[14]
    PIN A_DIN[18]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  266.97 0 267.23 0.26 ;
        END
    END A_DIN[18]
    PIN A_DIN[13]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  149.41 0 149.67 0.26 ;
        END
    END A_DIN[13]
    PIN A_BIST_DIN[18]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  266.115 0 266.375 0.26 ;
        END
    END A_BIST_DIN[18]
    PIN A_BIST_DIN[13]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  150.265 0 150.525 0.26 ;
        END
    END A_BIST_DIN[13]
    PIN A_BM[18]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  259.13 0 259.39 0.26 ;
        END
    END A_BM[18]
    PIN A_BM[13]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  157.25 0 157.51 0.26 ;
        END
    END A_BM[13]
    PIN A_BIST_BM[18]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  260.505 0 260.765 0.26 ;
        END
    END A_BIST_BM[18]
    PIN A_BIST_BM[13]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  155.875 0 156.135 0.26 ;
        END
    END A_BIST_BM[13]
    PIN A_DOUT[18]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  259.64 0 259.9 0.26 ;
        END
    END A_DOUT[18]
    PIN A_DOUT[13]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  156.74 0 157 0.26 ;
        END
    END A_DOUT[13]
    PIN A_DIN[19]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  278.21 0 278.47 0.26 ;
        END
    END A_DIN[19]
    PIN A_DIN[12]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  138.17 0 138.43 0.26 ;
        END
    END A_DIN[12]
    PIN A_BIST_DIN[19]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  277.355 0 277.615 0.26 ;
        END
    END A_BIST_DIN[19]
    PIN A_BIST_DIN[12]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  139.025 0 139.285 0.26 ;
        END
    END A_BIST_DIN[12]
    PIN A_BM[19]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  270.37 0 270.63 0.26 ;
        END
    END A_BM[19]
    PIN A_BM[12]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  146.01 0 146.27 0.26 ;
        END
    END A_BM[12]
    PIN A_BIST_BM[19]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  271.745 0 272.005 0.26 ;
        END
    END A_BIST_BM[19]
    PIN A_BIST_BM[12]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  144.635 0 144.895 0.26 ;
        END
    END A_BIST_BM[12]
    PIN A_DOUT[19]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  270.88 0 271.14 0.26 ;
        END
    END A_DOUT[19]
    PIN A_DOUT[12]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  145.5 0 145.76 0.26 ;
        END
    END A_DOUT[12]
    PIN A_DIN[20]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  289.45 0 289.71 0.26 ;
        END
    END A_DIN[20]
    PIN A_DIN[11]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  126.93 0 127.19 0.26 ;
        END
    END A_DIN[11]
    PIN A_BIST_DIN[20]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  288.595 0 288.855 0.26 ;
        END
    END A_BIST_DIN[20]
    PIN A_BIST_DIN[11]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  127.785 0 128.045 0.26 ;
        END
    END A_BIST_DIN[11]
    PIN A_BM[20]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  281.61 0 281.87 0.26 ;
        END
    END A_BM[20]
    PIN A_BM[11]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  134.77 0 135.03 0.26 ;
        END
    END A_BM[11]
    PIN A_BIST_BM[20]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  282.985 0 283.245 0.26 ;
        END
    END A_BIST_BM[20]
    PIN A_BIST_BM[11]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  133.395 0 133.655 0.26 ;
        END
    END A_BIST_BM[11]
    PIN A_DOUT[20]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  282.12 0 282.38 0.26 ;
        END
    END A_DOUT[20]
    PIN A_DOUT[11]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  134.26 0 134.52 0.26 ;
        END
    END A_DOUT[11]
    PIN A_DIN[21]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  300.69 0 300.95 0.26 ;
        END
    END A_DIN[21]
    PIN A_DIN[10]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  115.69 0 115.95 0.26 ;
        END
    END A_DIN[10]
    PIN A_BIST_DIN[21]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  299.835 0 300.095 0.26 ;
        END
    END A_BIST_DIN[21]
    PIN A_BIST_DIN[10]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  116.545 0 116.805 0.26 ;
        END
    END A_BIST_DIN[10]
    PIN A_BM[21]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  292.85 0 293.11 0.26 ;
        END
    END A_BM[21]
    PIN A_BM[10]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  123.53 0 123.79 0.26 ;
        END
    END A_BM[10]
    PIN A_BIST_BM[21]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  294.225 0 294.485 0.26 ;
        END
    END A_BIST_BM[21]
    PIN A_BIST_BM[10]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  122.155 0 122.415 0.26 ;
        END
    END A_BIST_BM[10]
    PIN A_DOUT[21]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  293.36 0 293.62 0.26 ;
        END
    END A_DOUT[21]
    PIN A_DOUT[10]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  123.02 0 123.28 0.26 ;
        END
    END A_DOUT[10]
    PIN A_DIN[22]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  311.93 0 312.19 0.26 ;
        END
    END A_DIN[22]
    PIN A_DIN[9]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  104.45 0 104.71 0.26 ;
        END
    END A_DIN[9]
    PIN A_BIST_DIN[22]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  311.075 0 311.335 0.26 ;
        END
    END A_BIST_DIN[22]
    PIN A_BIST_DIN[9]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  105.305 0 105.565 0.26 ;
        END
    END A_BIST_DIN[9]
    PIN A_BM[22]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  304.09 0 304.35 0.26 ;
        END
    END A_BM[22]
    PIN A_BM[9]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  112.29 0 112.55 0.26 ;
        END
    END A_BM[9]
    PIN A_BIST_BM[22]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  305.465 0 305.725 0.26 ;
        END
    END A_BIST_BM[22]
    PIN A_BIST_BM[9]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  110.915 0 111.175 0.26 ;
        END
    END A_BIST_BM[9]
    PIN A_DOUT[22]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  304.6 0 304.86 0.26 ;
        END
    END A_DOUT[22]
    PIN A_DOUT[9]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  111.78 0 112.04 0.26 ;
        END
    END A_DOUT[9]
    PIN A_DIN[23]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  323.17 0 323.43 0.26 ;
        END
    END A_DIN[23]
    PIN A_DIN[8]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  93.21 0 93.47 0.26 ;
        END
    END A_DIN[8]
    PIN A_BIST_DIN[23]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  322.315 0 322.575 0.26 ;
        END
    END A_BIST_DIN[23]
    PIN A_BIST_DIN[8]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  94.065 0 94.325 0.26 ;
        END
    END A_BIST_DIN[8]
    PIN A_BM[23]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  315.33 0 315.59 0.26 ;
        END
    END A_BM[23]
    PIN A_BM[8]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  101.05 0 101.31 0.26 ;
        END
    END A_BM[8]
    PIN A_BIST_BM[23]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  316.705 0 316.965 0.26 ;
        END
    END A_BIST_BM[23]
    PIN A_BIST_BM[8]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  99.675 0 99.935 0.26 ;
        END
    END A_BIST_BM[8]
    PIN A_DOUT[23]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  315.84 0 316.1 0.26 ;
        END
    END A_DOUT[23]
    PIN A_DOUT[8]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  100.54 0 100.8 0.26 ;
        END
    END A_DOUT[8]
    PIN A_DIN[24]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  334.41 0 334.67 0.26 ;
        END
    END A_DIN[24]
    PIN A_DIN[7]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  81.97 0 82.23 0.26 ;
        END
    END A_DIN[7]
    PIN A_BIST_DIN[24]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  333.555 0 333.815 0.26 ;
        END
    END A_BIST_DIN[24]
    PIN A_BIST_DIN[7]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  82.825 0 83.085 0.26 ;
        END
    END A_BIST_DIN[7]
    PIN A_BM[24]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  326.57 0 326.83 0.26 ;
        END
    END A_BM[24]
    PIN A_BM[7]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  89.81 0 90.07 0.26 ;
        END
    END A_BM[7]
    PIN A_BIST_BM[24]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  327.945 0 328.205 0.26 ;
        END
    END A_BIST_BM[24]
    PIN A_BIST_BM[7]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  88.435 0 88.695 0.26 ;
        END
    END A_BIST_BM[7]
    PIN A_DOUT[24]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  327.08 0 327.34 0.26 ;
        END
    END A_DOUT[24]
    PIN A_DOUT[7]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  89.3 0 89.56 0.26 ;
        END
    END A_DOUT[7]
    PIN A_DIN[25]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  345.65 0 345.91 0.26 ;
        END
    END A_DIN[25]
    PIN A_DIN[6]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  70.73 0 70.99 0.26 ;
        END
    END A_DIN[6]
    PIN A_BIST_DIN[25]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  344.795 0 345.055 0.26 ;
        END
    END A_BIST_DIN[25]
    PIN A_BIST_DIN[6]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  71.585 0 71.845 0.26 ;
        END
    END A_BIST_DIN[6]
    PIN A_BM[25]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  337.81 0 338.07 0.26 ;
        END
    END A_BM[25]
    PIN A_BM[6]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  78.57 0 78.83 0.26 ;
        END
    END A_BM[6]
    PIN A_BIST_BM[25]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  339.185 0 339.445 0.26 ;
        END
    END A_BIST_BM[25]
    PIN A_BIST_BM[6]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  77.195 0 77.455 0.26 ;
        END
    END A_BIST_BM[6]
    PIN A_DOUT[25]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  338.32 0 338.58 0.26 ;
        END
    END A_DOUT[25]
    PIN A_DOUT[6]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  78.06 0 78.32 0.26 ;
        END
    END A_DOUT[6]
    PIN A_DIN[26]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  356.89 0 357.15 0.26 ;
        END
    END A_DIN[26]
    PIN A_DIN[5]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  59.49 0 59.75 0.26 ;
        END
    END A_DIN[5]
    PIN A_BIST_DIN[26]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  356.035 0 356.295 0.26 ;
        END
    END A_BIST_DIN[26]
    PIN A_BIST_DIN[5]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  60.345 0 60.605 0.26 ;
        END
    END A_BIST_DIN[5]
    PIN A_BM[26]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  349.05 0 349.31 0.26 ;
        END
    END A_BM[26]
    PIN A_BM[5]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  67.33 0 67.59 0.26 ;
        END
    END A_BM[5]
    PIN A_BIST_BM[26]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  350.425 0 350.685 0.26 ;
        END
    END A_BIST_BM[26]
    PIN A_BIST_BM[5]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  65.955 0 66.215 0.26 ;
        END
    END A_BIST_BM[5]
    PIN A_DOUT[26]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  349.56 0 349.82 0.26 ;
        END
    END A_DOUT[26]
    PIN A_DOUT[5]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  66.82 0 67.08 0.26 ;
        END
    END A_DOUT[5]
    PIN A_DIN[27]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  368.13 0 368.39 0.26 ;
        END
    END A_DIN[27]
    PIN A_DIN[4]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  48.25 0 48.51 0.26 ;
        END
    END A_DIN[4]
    PIN A_BIST_DIN[27]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  367.275 0 367.535 0.26 ;
        END
    END A_BIST_DIN[27]
    PIN A_BIST_DIN[4]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  49.105 0 49.365 0.26 ;
        END
    END A_BIST_DIN[4]
    PIN A_BM[27]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  360.29 0 360.55 0.26 ;
        END
    END A_BM[27]
    PIN A_BM[4]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  56.09 0 56.35 0.26 ;
        END
    END A_BM[4]
    PIN A_BIST_BM[27]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  361.665 0 361.925 0.26 ;
        END
    END A_BIST_BM[27]
    PIN A_BIST_BM[4]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  54.715 0 54.975 0.26 ;
        END
    END A_BIST_BM[4]
    PIN A_DOUT[27]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  360.8 0 361.06 0.26 ;
        END
    END A_DOUT[27]
    PIN A_DOUT[4]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  55.58 0 55.84 0.26 ;
        END
    END A_DOUT[4]
    PIN A_DIN[28]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  379.37 0 379.63 0.26 ;
        END
    END A_DIN[28]
    PIN A_DIN[3]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  37.01 0 37.27 0.26 ;
        END
    END A_DIN[3]
    PIN A_BIST_DIN[28]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  378.515 0 378.775 0.26 ;
        END
    END A_BIST_DIN[28]
    PIN A_BIST_DIN[3]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  37.865 0 38.125 0.26 ;
        END
    END A_BIST_DIN[3]
    PIN A_BM[28]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  371.53 0 371.79 0.26 ;
        END
    END A_BM[28]
    PIN A_BM[3]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  44.85 0 45.11 0.26 ;
        END
    END A_BM[3]
    PIN A_BIST_BM[28]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  372.905 0 373.165 0.26 ;
        END
    END A_BIST_BM[28]
    PIN A_BIST_BM[3]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  43.475 0 43.735 0.26 ;
        END
    END A_BIST_BM[3]
    PIN A_DOUT[28]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  372.04 0 372.3 0.26 ;
        END
    END A_DOUT[28]
    PIN A_DOUT[3]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  44.34 0 44.6 0.26 ;
        END
    END A_DOUT[3]
    PIN A_DIN[29]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  390.61 0 390.87 0.26 ;
        END
    END A_DIN[29]
    PIN A_DIN[2]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  25.77 0 26.03 0.26 ;
        END
    END A_DIN[2]
    PIN A_BIST_DIN[29]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  389.755 0 390.015 0.26 ;
        END
    END A_BIST_DIN[29]
    PIN A_BIST_DIN[2]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  26.625 0 26.885 0.26 ;
        END
    END A_BIST_DIN[2]
    PIN A_BM[29]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  382.77 0 383.03 0.26 ;
        END
    END A_BM[29]
    PIN A_BM[2]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  33.61 0 33.87 0.26 ;
        END
    END A_BM[2]
    PIN A_BIST_BM[29]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  384.145 0 384.405 0.26 ;
        END
    END A_BIST_BM[29]
    PIN A_BIST_BM[2]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  32.235 0 32.495 0.26 ;
        END
    END A_BIST_BM[2]
    PIN A_DOUT[29]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  383.28 0 383.54 0.26 ;
        END
    END A_DOUT[29]
    PIN A_DOUT[2]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  33.1 0 33.36 0.26 ;
        END
    END A_DOUT[2]
    PIN A_DIN[30]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  401.85 0 402.11 0.26 ;
        END
    END A_DIN[30]
    PIN A_DIN[1]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  14.53 0 14.79 0.26 ;
        END
    END A_DIN[1]
    PIN A_BIST_DIN[30]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  400.995 0 401.255 0.26 ;
        END
    END A_BIST_DIN[30]
    PIN A_BIST_DIN[1]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  15.385 0 15.645 0.26 ;
        END
    END A_BIST_DIN[1]
    PIN A_BM[30]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  394.01 0 394.27 0.26 ;
        END
    END A_BM[30]
    PIN A_BM[1]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  22.37 0 22.63 0.26 ;
        END
    END A_BM[1]
    PIN A_BIST_BM[30]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  395.385 0 395.645 0.26 ;
        END
    END A_BIST_BM[30]
    PIN A_BIST_BM[1]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  20.995 0 21.255 0.26 ;
        END
    END A_BIST_BM[1]
    PIN A_DOUT[30]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  394.52 0 394.78 0.26 ;
        END
    END A_DOUT[30]
    PIN A_DOUT[1]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  21.86 0 22.12 0.26 ;
        END
    END A_DOUT[1]
    PIN A_DIN[31]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  413.09 0 413.35 0.26 ;
        END
    END A_DIN[31]
    PIN A_DIN[0]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  3.29 0 3.55 0.26 ;
        END
    END A_DIN[0]
    PIN A_BIST_DIN[31]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  412.235 0 412.495 0.26 ;
        END
    END A_BIST_DIN[31]
    PIN A_BIST_DIN[0]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  4.145 0 4.405 0.26 ;
        END
    END A_BIST_DIN[0]
    PIN A_BM[31]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  405.25 0 405.51 0.26 ;
        END
    END A_BM[31]
    PIN A_BM[0]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  11.13 0 11.39 0.26 ;
        END
    END A_BM[0]
    PIN A_BIST_BM[31]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  406.625 0 406.885 0.26 ;
        END
    END A_BIST_BM[31]
    PIN A_BIST_BM[0]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  9.755 0 10.015 0.26 ;
        END
    END A_BIST_BM[0]
    PIN A_DOUT[31]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  405.76 0 406.02 0.26 ;
        END
    END A_DOUT[31]
    PIN A_DOUT[0]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  10.62 0 10.88 0.26 ;
        END
    END A_DOUT[0]
    PIN A_ADDR[0]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 8.9011 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 45.2233 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  204.52 0 204.78 0.26 ;
        END
    END A_ADDR[0]
    PIN A_BIST_ADDR[0]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 9.6967 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 49.1845 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  209.11 0 209.37 0.26 ;
        END
    END A_BIST_ADDR[0]
    PIN A_ADDR[1]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 7.774 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 39.657 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  204.01 0 204.27 0.26 ;
        END
    END A_ADDR[1]
    PIN A_BIST_ADDR[1]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 8.5696 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 43.6181 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  208.6 0 208.86 0.26 ;
        END
    END A_BIST_ADDR[1]
    PIN A_ADDR[2]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 10.6327 LAYER Metal2 ;
        ANTENNAPARTIALMETALAREA 1.5246 LAYER Metal3 ;
        ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
        ANTENNAMAXAREACAR 9.41598 LAYER Metal3 ;
        PORT
            LAYER Metal2 ;
              RECT  212.17 0 212.43 0.26 ;
        END
    END A_ADDR[2]
    PIN A_BIST_ADDR[2]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 10.6327 LAYER Metal2 ;
        ANTENNAPARTIALMETALAREA 1.0962 LAYER Metal3 ;
        ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
        ANTENNAMAXAREACAR 7.81379 LAYER Metal3 ;
        PORT
            LAYER Metal2 ;
              RECT  212.68 0 212.94 0.26 ;
        END
    END A_BIST_ADDR[2]
    PIN A_ADDR[3]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 10.6327 LAYER Metal2 ;
        ANTENNAPARTIALMETALAREA 3.8367 LAYER Metal3 ;
        ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
        ANTENNAMAXAREACAR 20.9276 LAYER Metal3 ;
        PORT
            LAYER Metal2 ;
              RECT  211.15 0 211.41 0.26 ;
        END
    END A_ADDR[3]
    PIN A_BIST_ADDR[3]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 10.6327 LAYER Metal2 ;
        ANTENNAPARTIALMETALAREA 3.5175 LAYER Metal3 ;
        ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
        ANTENNAMAXAREACAR 19.8691 LAYER Metal3 ;
        PORT
            LAYER Metal2 ;
              RECT  211.66 0 211.92 0.26 ;
        END
    END A_BIST_ADDR[3]
    PIN A_ADDR[4]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 12.1979 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 61.6375 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  214.72 0 214.98 0.26 ;
        END
    END A_ADDR[4]
    PIN A_BIST_ADDR[4]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 11.9327 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 60.3172 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  214.21 0 214.47 0.26 ;
        END
    END A_BIST_ADDR[4]
    PIN A_ADDR[5]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 13.9269 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 70.246 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  213.7 0 213.96 0.26 ;
        END
    END A_ADDR[5]
    PIN A_BIST_ADDR[5]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 13.6617 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 68.9256 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  213.19 0 213.45 0.26 ;
        END
    END A_BIST_ADDR[5]
    PIN A_ADDR[6]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 10.9525 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 55.4369 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  192.28 0 192.54 0.26 ;
        END
    END A_ADDR[6]
    PIN A_BIST_ADDR[6]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 10.6771 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 54.0657 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  192.79 0 193.05 0.26 ;
        END
    END A_BIST_ADDR[6]
    PIN A_ADDR[7]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 12.4163 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 62.7249 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  193.3 0 193.56 0.26 ;
        END
    END A_ADDR[7]
    PIN A_BIST_ADDR[7]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 12.1511 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 61.4045 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  193.81 0 194.07 0.26 ;
        END
    END A_BIST_ADDR[7]
    PIN A_ADDR[8]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 10.3675 LAYER Metal2 ;
        ANTENNAPARTIALMETALAREA 1.5897 LAYER Metal3 ;
        ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
        ANTENNAMAXAREACAR 9.7401 LAYER Metal3 ;
        PORT
            LAYER Metal2 ;
              RECT  222.37 0 222.63 0.26 ;
        END
    END A_ADDR[8]
    PIN A_BIST_ADDR[8]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 10.3675 LAYER Metal2 ;
        ANTENNAPARTIALMETALAREA 1.3755 LAYER Metal3 ;
        ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
        ANTENNAMAXAREACAR 9.20438 LAYER Metal3 ;
        PORT
            LAYER Metal2 ;
              RECT  222.88 0 223.14 0.26 ;
        END
    END A_BIST_ADDR[8]
    PIN A_CLK
        DIRECTION INPUT ; 
        USE CLOCK ; 
        ANTENNAPARTIALMETALAREA 4.0547 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 21.0939 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  202.48 0 202.74 0.26 ;
        END
    END A_CLK
    PIN A_REN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.99505 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 20.7969 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  206.05 0 206.31 0.26 ;
        END
    END A_REN
    PIN A_WEN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 15.2686 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  205.54 0 205.8 0.26 ;
        END
    END A_WEN
    PIN A_MEN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.0247 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 15.9656 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  202.99 0 203.25 0.26 ;
        END
    END A_MEN
    PIN A_DLY
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 6.058 LAYER Metal2 ;
        ANTENNAGATEAREA 0.3367 LAYER Metal2 ;
        ANTENNAMAXAREACAR 18.5328 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  224.41 0 224.67 0.26 ;
        END
    END A_DLY
    PIN A_BIST_EN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.9871 LAYER Metal2 ;
        ANTENNAPARTIALMETALAREA 203.317 LAYER Metal3 ;
        ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
        ANTENNAGATEAREA 1.43 LAYER Metal2 ;
        ANTENNAGATEAREA 27.5275 LAYER Metal3 ;
        ANTENNAMAXAREACAR 3.21364 LAYER Metal2 ;
        ANTENNAMAXAREACAR 17.6587 LAYER Metal3 ;
        ANTENNAMAXCUTCAR 0.151469 LAYER Via2 ;
        PORT
            LAYER Metal2 ;
              RECT  205.03 0 205.29 0.26 ;
        END
    END A_BIST_EN
    PIN A_BIST_CLK
        DIRECTION INPUT ; 
        USE CLOCK ; 
        ANTENNAPARTIALMETALAREA 4.1639 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 21.9534 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  200.95 0 201.21 0.26 ;
        END
    END A_BIST_CLK
    PIN A_BIST_REN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 4.1119 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 21.6945 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  207.58 0 207.84 0.26 ;
        END
    END A_BIST_REN
    PIN A_BIST_WEN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 2.9051 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 15.6861 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  207.07 0 207.33 0.26 ;
        END
    END A_BIST_WEN
    PIN A_BIST_MEN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 2.8977 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 15.6492 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  201.46 0 201.72 0.26 ;
        END
    END A_BIST_MEN
    OBS
      LAYER Metal1 ;
        RECT  0 0 416.64 191.34 ;
      LAYER Metal2 ;
        RECT  0.105 45.465 0.305 191.315 ;
        RECT  1.1 190.585 1.3 191.315 ;
        RECT  3.29 0.52 3.55 5.16 ;
        RECT  2.77 4.9 3.55 5.16 ;
        RECT  2.77 4.9 3.03 6.64 ;
        RECT  1.92 190.585 2.12 191.315 ;
        RECT  2.415 190.585 2.615 191.315 ;
        RECT  2.915 190.585 3.115 191.315 ;
        RECT  3.415 190.585 3.615 191.315 ;
        RECT  3.91 190.585 4.11 191.315 ;
        RECT  4.655 0.17 5.425 0.94 ;
        RECT  4.655 0.17 4.915 12.9 ;
        RECT  5.165 0.17 5.425 12.9 ;
        RECT  4.145 0.52 4.405 5.815 ;
        RECT  4.73 190.585 4.93 191.315 ;
        RECT  5.675 0.17 6.445 0.43 ;
        RECT  5.675 0.17 5.935 11.5 ;
        RECT  6.185 0.17 6.445 11.5 ;
        RECT  5.225 190.585 5.425 191.315 ;
        RECT  5.725 190.585 5.925 191.315 ;
        RECT  6.225 190.585 6.425 191.315 ;
        RECT  7.715 0.17 8.485 0.43 ;
        RECT  7.715 0.17 7.975 10.48 ;
        RECT  8.225 0.17 8.485 10.99 ;
        RECT  6.72 190.585 6.92 191.315 ;
        RECT  7.54 190.585 7.74 191.315 ;
        RECT  8.735 0.17 9.505 0.94 ;
        RECT  8.735 0.17 8.995 8.7 ;
        RECT  9.245 0.17 9.505 12.9 ;
        RECT  8.035 190.585 8.235 191.315 ;
        RECT  8.535 190.585 8.735 191.315 ;
        RECT  9.035 190.585 9.235 191.315 ;
        RECT  9.53 190.585 9.73 191.315 ;
        RECT  9.755 0.52 10.015 2.485 ;
        RECT  10.35 190.585 10.55 191.315 ;
        RECT  10.62 0.52 10.88 14.11 ;
        RECT  10.845 190.585 11.045 191.315 ;
        RECT  11.13 0.52 11.39 2.335 ;
        RECT  11.345 190.585 11.545 191.315 ;
        RECT  11.845 190.585 12.045 191.315 ;
        RECT  12.34 190.585 12.54 191.315 ;
        RECT  14.53 0.52 14.79 5.16 ;
        RECT  14.01 4.9 14.79 5.16 ;
        RECT  14.01 4.9 14.27 6.64 ;
        RECT  13.16 190.585 13.36 191.315 ;
        RECT  13.655 190.585 13.855 191.315 ;
        RECT  14.155 190.585 14.355 191.315 ;
        RECT  14.655 190.585 14.855 191.315 ;
        RECT  15.15 190.585 15.35 191.315 ;
        RECT  15.895 0.17 16.665 0.94 ;
        RECT  15.895 0.17 16.155 12.9 ;
        RECT  16.405 0.17 16.665 12.9 ;
        RECT  15.385 0.52 15.645 5.815 ;
        RECT  15.97 190.585 16.17 191.315 ;
        RECT  16.915 0.17 17.685 0.43 ;
        RECT  16.915 0.17 17.175 11.5 ;
        RECT  17.425 0.17 17.685 11.5 ;
        RECT  16.465 190.585 16.665 191.315 ;
        RECT  16.965 190.585 17.165 191.315 ;
        RECT  17.465 190.585 17.665 191.315 ;
        RECT  18.955 0.17 19.725 0.43 ;
        RECT  18.955 0.17 19.215 10.48 ;
        RECT  19.465 0.17 19.725 10.99 ;
        RECT  17.96 190.585 18.16 191.315 ;
        RECT  18.78 190.585 18.98 191.315 ;
        RECT  19.975 0.17 20.745 0.94 ;
        RECT  19.975 0.17 20.235 8.7 ;
        RECT  20.485 0.17 20.745 12.9 ;
        RECT  19.275 190.585 19.475 191.315 ;
        RECT  19.775 190.585 19.975 191.315 ;
        RECT  20.275 190.585 20.475 191.315 ;
        RECT  20.77 190.585 20.97 191.315 ;
        RECT  20.995 0.52 21.255 2.485 ;
        RECT  21.59 190.585 21.79 191.315 ;
        RECT  21.86 0.52 22.12 14.11 ;
        RECT  22.085 190.585 22.285 191.315 ;
        RECT  22.37 0.52 22.63 2.335 ;
        RECT  22.585 190.585 22.785 191.315 ;
        RECT  23.085 190.585 23.285 191.315 ;
        RECT  23.58 190.585 23.78 191.315 ;
        RECT  25.77 0.52 26.03 5.16 ;
        RECT  25.25 4.9 26.03 5.16 ;
        RECT  25.25 4.9 25.51 6.64 ;
        RECT  24.4 190.585 24.6 191.315 ;
        RECT  24.895 190.585 25.095 191.315 ;
        RECT  25.395 190.585 25.595 191.315 ;
        RECT  25.895 190.585 26.095 191.315 ;
        RECT  26.39 190.585 26.59 191.315 ;
        RECT  27.135 0.17 27.905 0.94 ;
        RECT  27.135 0.17 27.395 12.9 ;
        RECT  27.645 0.17 27.905 12.9 ;
        RECT  26.625 0.52 26.885 5.815 ;
        RECT  27.21 190.585 27.41 191.315 ;
        RECT  28.155 0.17 28.925 0.43 ;
        RECT  28.155 0.17 28.415 11.5 ;
        RECT  28.665 0.17 28.925 11.5 ;
        RECT  27.705 190.585 27.905 191.315 ;
        RECT  28.205 190.585 28.405 191.315 ;
        RECT  28.705 190.585 28.905 191.315 ;
        RECT  30.195 0.17 30.965 0.43 ;
        RECT  30.195 0.17 30.455 10.48 ;
        RECT  30.705 0.17 30.965 10.99 ;
        RECT  29.2 190.585 29.4 191.315 ;
        RECT  30.02 190.585 30.22 191.315 ;
        RECT  31.215 0.17 31.985 0.94 ;
        RECT  31.215 0.17 31.475 8.7 ;
        RECT  31.725 0.17 31.985 12.9 ;
        RECT  30.515 190.585 30.715 191.315 ;
        RECT  31.015 190.585 31.215 191.315 ;
        RECT  31.515 190.585 31.715 191.315 ;
        RECT  32.01 190.585 32.21 191.315 ;
        RECT  32.235 0.52 32.495 2.485 ;
        RECT  32.83 190.585 33.03 191.315 ;
        RECT  33.1 0.52 33.36 14.11 ;
        RECT  33.325 190.585 33.525 191.315 ;
        RECT  33.61 0.52 33.87 2.335 ;
        RECT  33.825 190.585 34.025 191.315 ;
        RECT  34.325 190.585 34.525 191.315 ;
        RECT  34.82 190.585 35.02 191.315 ;
        RECT  37.01 0.52 37.27 5.16 ;
        RECT  36.49 4.9 37.27 5.16 ;
        RECT  36.49 4.9 36.75 6.64 ;
        RECT  35.64 190.585 35.84 191.315 ;
        RECT  36.135 190.585 36.335 191.315 ;
        RECT  36.635 190.585 36.835 191.315 ;
        RECT  37.135 190.585 37.335 191.315 ;
        RECT  37.63 190.585 37.83 191.315 ;
        RECT  38.375 0.17 39.145 0.94 ;
        RECT  38.375 0.17 38.635 12.9 ;
        RECT  38.885 0.17 39.145 12.9 ;
        RECT  37.865 0.52 38.125 5.815 ;
        RECT  38.45 190.585 38.65 191.315 ;
        RECT  39.395 0.17 40.165 0.43 ;
        RECT  39.395 0.17 39.655 11.5 ;
        RECT  39.905 0.17 40.165 11.5 ;
        RECT  38.945 190.585 39.145 191.315 ;
        RECT  39.445 190.585 39.645 191.315 ;
        RECT  39.945 190.585 40.145 191.315 ;
        RECT  41.435 0.17 42.205 0.43 ;
        RECT  41.435 0.17 41.695 10.48 ;
        RECT  41.945 0.17 42.205 10.99 ;
        RECT  40.44 190.585 40.64 191.315 ;
        RECT  41.26 190.585 41.46 191.315 ;
        RECT  42.455 0.17 43.225 0.94 ;
        RECT  42.455 0.17 42.715 8.7 ;
        RECT  42.965 0.17 43.225 12.9 ;
        RECT  41.755 190.585 41.955 191.315 ;
        RECT  42.255 190.585 42.455 191.315 ;
        RECT  42.755 190.585 42.955 191.315 ;
        RECT  43.25 190.585 43.45 191.315 ;
        RECT  43.475 0.52 43.735 2.485 ;
        RECT  44.07 190.585 44.27 191.315 ;
        RECT  44.34 0.52 44.6 14.11 ;
        RECT  44.565 190.585 44.765 191.315 ;
        RECT  44.85 0.52 45.11 2.335 ;
        RECT  45.065 190.585 45.265 191.315 ;
        RECT  45.565 190.585 45.765 191.315 ;
        RECT  46.06 190.585 46.26 191.315 ;
        RECT  48.25 0.52 48.51 5.16 ;
        RECT  47.73 4.9 48.51 5.16 ;
        RECT  47.73 4.9 47.99 6.64 ;
        RECT  46.88 190.585 47.08 191.315 ;
        RECT  47.375 190.585 47.575 191.315 ;
        RECT  47.875 190.585 48.075 191.315 ;
        RECT  48.375 190.585 48.575 191.315 ;
        RECT  48.87 190.585 49.07 191.315 ;
        RECT  49.615 0.17 50.385 0.94 ;
        RECT  49.615 0.17 49.875 12.9 ;
        RECT  50.125 0.17 50.385 12.9 ;
        RECT  49.105 0.52 49.365 5.815 ;
        RECT  49.69 190.585 49.89 191.315 ;
        RECT  50.635 0.17 51.405 0.43 ;
        RECT  50.635 0.17 50.895 11.5 ;
        RECT  51.145 0.17 51.405 11.5 ;
        RECT  50.185 190.585 50.385 191.315 ;
        RECT  50.685 190.585 50.885 191.315 ;
        RECT  51.185 190.585 51.385 191.315 ;
        RECT  52.675 0.17 53.445 0.43 ;
        RECT  52.675 0.17 52.935 10.48 ;
        RECT  53.185 0.17 53.445 10.99 ;
        RECT  51.68 190.585 51.88 191.315 ;
        RECT  52.5 190.585 52.7 191.315 ;
        RECT  53.695 0.17 54.465 0.94 ;
        RECT  53.695 0.17 53.955 8.7 ;
        RECT  54.205 0.17 54.465 12.9 ;
        RECT  52.995 190.585 53.195 191.315 ;
        RECT  53.495 190.585 53.695 191.315 ;
        RECT  53.995 190.585 54.195 191.315 ;
        RECT  54.49 190.585 54.69 191.315 ;
        RECT  54.715 0.52 54.975 2.485 ;
        RECT  55.31 190.585 55.51 191.315 ;
        RECT  55.58 0.52 55.84 14.11 ;
        RECT  55.805 190.585 56.005 191.315 ;
        RECT  56.09 0.52 56.35 2.335 ;
        RECT  56.305 190.585 56.505 191.315 ;
        RECT  56.805 190.585 57.005 191.315 ;
        RECT  57.3 190.585 57.5 191.315 ;
        RECT  59.49 0.52 59.75 5.16 ;
        RECT  58.97 4.9 59.75 5.16 ;
        RECT  58.97 4.9 59.23 6.64 ;
        RECT  58.12 190.585 58.32 191.315 ;
        RECT  58.615 190.585 58.815 191.315 ;
        RECT  59.115 190.585 59.315 191.315 ;
        RECT  59.615 190.585 59.815 191.315 ;
        RECT  60.11 190.585 60.31 191.315 ;
        RECT  60.855 0.17 61.625 0.94 ;
        RECT  60.855 0.17 61.115 12.9 ;
        RECT  61.365 0.17 61.625 12.9 ;
        RECT  60.345 0.52 60.605 5.815 ;
        RECT  60.93 190.585 61.13 191.315 ;
        RECT  61.875 0.17 62.645 0.43 ;
        RECT  61.875 0.17 62.135 11.5 ;
        RECT  62.385 0.17 62.645 11.5 ;
        RECT  61.425 190.585 61.625 191.315 ;
        RECT  61.925 190.585 62.125 191.315 ;
        RECT  62.425 190.585 62.625 191.315 ;
        RECT  63.915 0.17 64.685 0.43 ;
        RECT  63.915 0.17 64.175 10.48 ;
        RECT  64.425 0.17 64.685 10.99 ;
        RECT  62.92 190.585 63.12 191.315 ;
        RECT  63.74 190.585 63.94 191.315 ;
        RECT  64.935 0.17 65.705 0.94 ;
        RECT  64.935 0.17 65.195 8.7 ;
        RECT  65.445 0.17 65.705 12.9 ;
        RECT  64.235 190.585 64.435 191.315 ;
        RECT  64.735 190.585 64.935 191.315 ;
        RECT  65.235 190.585 65.435 191.315 ;
        RECT  65.73 190.585 65.93 191.315 ;
        RECT  65.955 0.52 66.215 2.485 ;
        RECT  66.55 190.585 66.75 191.315 ;
        RECT  66.82 0.52 67.08 14.11 ;
        RECT  67.045 190.585 67.245 191.315 ;
        RECT  67.33 0.52 67.59 2.335 ;
        RECT  67.545 190.585 67.745 191.315 ;
        RECT  68.045 190.585 68.245 191.315 ;
        RECT  68.54 190.585 68.74 191.315 ;
        RECT  70.73 0.52 70.99 5.16 ;
        RECT  70.21 4.9 70.99 5.16 ;
        RECT  70.21 4.9 70.47 6.64 ;
        RECT  69.36 190.585 69.56 191.315 ;
        RECT  69.855 190.585 70.055 191.315 ;
        RECT  70.355 190.585 70.555 191.315 ;
        RECT  70.855 190.585 71.055 191.315 ;
        RECT  71.35 190.585 71.55 191.315 ;
        RECT  72.095 0.17 72.865 0.94 ;
        RECT  72.095 0.17 72.355 12.9 ;
        RECT  72.605 0.17 72.865 12.9 ;
        RECT  71.585 0.52 71.845 5.815 ;
        RECT  72.17 190.585 72.37 191.315 ;
        RECT  73.115 0.17 73.885 0.43 ;
        RECT  73.115 0.17 73.375 11.5 ;
        RECT  73.625 0.17 73.885 11.5 ;
        RECT  72.665 190.585 72.865 191.315 ;
        RECT  73.165 190.585 73.365 191.315 ;
        RECT  73.665 190.585 73.865 191.315 ;
        RECT  75.155 0.17 75.925 0.43 ;
        RECT  75.155 0.17 75.415 10.48 ;
        RECT  75.665 0.17 75.925 10.99 ;
        RECT  74.16 190.585 74.36 191.315 ;
        RECT  74.98 190.585 75.18 191.315 ;
        RECT  76.175 0.17 76.945 0.94 ;
        RECT  76.175 0.17 76.435 8.7 ;
        RECT  76.685 0.17 76.945 12.9 ;
        RECT  75.475 190.585 75.675 191.315 ;
        RECT  75.975 190.585 76.175 191.315 ;
        RECT  76.475 190.585 76.675 191.315 ;
        RECT  76.97 190.585 77.17 191.315 ;
        RECT  77.195 0.52 77.455 2.485 ;
        RECT  77.79 190.585 77.99 191.315 ;
        RECT  78.06 0.52 78.32 14.11 ;
        RECT  78.285 190.585 78.485 191.315 ;
        RECT  78.57 0.52 78.83 2.335 ;
        RECT  78.785 190.585 78.985 191.315 ;
        RECT  79.285 190.585 79.485 191.315 ;
        RECT  79.78 190.585 79.98 191.315 ;
        RECT  81.97 0.52 82.23 5.16 ;
        RECT  81.45 4.9 82.23 5.16 ;
        RECT  81.45 4.9 81.71 6.64 ;
        RECT  80.6 190.585 80.8 191.315 ;
        RECT  81.095 190.585 81.295 191.315 ;
        RECT  81.595 190.585 81.795 191.315 ;
        RECT  82.095 190.585 82.295 191.315 ;
        RECT  82.59 190.585 82.79 191.315 ;
        RECT  83.335 0.17 84.105 0.94 ;
        RECT  83.335 0.17 83.595 12.9 ;
        RECT  83.845 0.17 84.105 12.9 ;
        RECT  82.825 0.52 83.085 5.815 ;
        RECT  83.41 190.585 83.61 191.315 ;
        RECT  84.355 0.17 85.125 0.43 ;
        RECT  84.355 0.17 84.615 11.5 ;
        RECT  84.865 0.17 85.125 11.5 ;
        RECT  83.905 190.585 84.105 191.315 ;
        RECT  84.405 190.585 84.605 191.315 ;
        RECT  84.905 190.585 85.105 191.315 ;
        RECT  86.395 0.17 87.165 0.43 ;
        RECT  86.395 0.17 86.655 10.48 ;
        RECT  86.905 0.17 87.165 10.99 ;
        RECT  85.4 190.585 85.6 191.315 ;
        RECT  86.22 190.585 86.42 191.315 ;
        RECT  87.415 0.17 88.185 0.94 ;
        RECT  87.415 0.17 87.675 8.7 ;
        RECT  87.925 0.17 88.185 12.9 ;
        RECT  86.715 190.585 86.915 191.315 ;
        RECT  87.215 190.585 87.415 191.315 ;
        RECT  87.715 190.585 87.915 191.315 ;
        RECT  88.21 190.585 88.41 191.315 ;
        RECT  88.435 0.52 88.695 2.485 ;
        RECT  89.03 190.585 89.23 191.315 ;
        RECT  89.3 0.52 89.56 14.11 ;
        RECT  89.525 190.585 89.725 191.315 ;
        RECT  89.81 0.52 90.07 2.335 ;
        RECT  90.025 190.585 90.225 191.315 ;
        RECT  90.525 190.585 90.725 191.315 ;
        RECT  91.02 190.585 91.22 191.315 ;
        RECT  93.21 0.52 93.47 5.16 ;
        RECT  92.69 4.9 93.47 5.16 ;
        RECT  92.69 4.9 92.95 6.64 ;
        RECT  91.84 190.585 92.04 191.315 ;
        RECT  92.335 190.585 92.535 191.315 ;
        RECT  92.835 190.585 93.035 191.315 ;
        RECT  93.335 190.585 93.535 191.315 ;
        RECT  93.83 190.585 94.03 191.315 ;
        RECT  94.575 0.17 95.345 0.94 ;
        RECT  94.575 0.17 94.835 12.9 ;
        RECT  95.085 0.17 95.345 12.9 ;
        RECT  94.065 0.52 94.325 5.815 ;
        RECT  94.65 190.585 94.85 191.315 ;
        RECT  95.595 0.17 96.365 0.43 ;
        RECT  95.595 0.17 95.855 11.5 ;
        RECT  96.105 0.17 96.365 11.5 ;
        RECT  95.145 190.585 95.345 191.315 ;
        RECT  95.645 190.585 95.845 191.315 ;
        RECT  96.145 190.585 96.345 191.315 ;
        RECT  97.635 0.17 98.405 0.43 ;
        RECT  97.635 0.17 97.895 10.48 ;
        RECT  98.145 0.17 98.405 10.99 ;
        RECT  96.64 190.585 96.84 191.315 ;
        RECT  97.46 190.585 97.66 191.315 ;
        RECT  98.655 0.17 99.425 0.94 ;
        RECT  98.655 0.17 98.915 8.7 ;
        RECT  99.165 0.17 99.425 12.9 ;
        RECT  97.955 190.585 98.155 191.315 ;
        RECT  98.455 190.585 98.655 191.315 ;
        RECT  98.955 190.585 99.155 191.315 ;
        RECT  99.45 190.585 99.65 191.315 ;
        RECT  99.675 0.52 99.935 2.485 ;
        RECT  100.27 190.585 100.47 191.315 ;
        RECT  100.54 0.52 100.8 14.11 ;
        RECT  100.765 190.585 100.965 191.315 ;
        RECT  101.05 0.52 101.31 2.335 ;
        RECT  101.265 190.585 101.465 191.315 ;
        RECT  101.765 190.585 101.965 191.315 ;
        RECT  102.26 190.585 102.46 191.315 ;
        RECT  104.45 0.52 104.71 5.16 ;
        RECT  103.93 4.9 104.71 5.16 ;
        RECT  103.93 4.9 104.19 6.64 ;
        RECT  103.08 190.585 103.28 191.315 ;
        RECT  103.575 190.585 103.775 191.315 ;
        RECT  104.075 190.585 104.275 191.315 ;
        RECT  104.575 190.585 104.775 191.315 ;
        RECT  105.07 190.585 105.27 191.315 ;
        RECT  105.815 0.17 106.585 0.94 ;
        RECT  105.815 0.17 106.075 12.9 ;
        RECT  106.325 0.17 106.585 12.9 ;
        RECT  105.305 0.52 105.565 5.815 ;
        RECT  105.89 190.585 106.09 191.315 ;
        RECT  106.835 0.17 107.605 0.43 ;
        RECT  106.835 0.17 107.095 11.5 ;
        RECT  107.345 0.17 107.605 11.5 ;
        RECT  106.385 190.585 106.585 191.315 ;
        RECT  106.885 190.585 107.085 191.315 ;
        RECT  107.385 190.585 107.585 191.315 ;
        RECT  108.875 0.17 109.645 0.43 ;
        RECT  108.875 0.17 109.135 10.48 ;
        RECT  109.385 0.17 109.645 10.99 ;
        RECT  107.88 190.585 108.08 191.315 ;
        RECT  108.7 190.585 108.9 191.315 ;
        RECT  109.895 0.17 110.665 0.94 ;
        RECT  109.895 0.17 110.155 8.7 ;
        RECT  110.405 0.17 110.665 12.9 ;
        RECT  109.195 190.585 109.395 191.315 ;
        RECT  109.695 190.585 109.895 191.315 ;
        RECT  110.195 190.585 110.395 191.315 ;
        RECT  110.69 190.585 110.89 191.315 ;
        RECT  110.915 0.52 111.175 2.485 ;
        RECT  111.51 190.585 111.71 191.315 ;
        RECT  111.78 0.52 112.04 14.11 ;
        RECT  112.005 190.585 112.205 191.315 ;
        RECT  112.29 0.52 112.55 2.335 ;
        RECT  112.505 190.585 112.705 191.315 ;
        RECT  113.005 190.585 113.205 191.315 ;
        RECT  113.5 190.585 113.7 191.315 ;
        RECT  115.69 0.52 115.95 5.16 ;
        RECT  115.17 4.9 115.95 5.16 ;
        RECT  115.17 4.9 115.43 6.64 ;
        RECT  114.32 190.585 114.52 191.315 ;
        RECT  114.815 190.585 115.015 191.315 ;
        RECT  115.315 190.585 115.515 191.315 ;
        RECT  115.815 190.585 116.015 191.315 ;
        RECT  116.31 190.585 116.51 191.315 ;
        RECT  117.055 0.17 117.825 0.94 ;
        RECT  117.055 0.17 117.315 12.9 ;
        RECT  117.565 0.17 117.825 12.9 ;
        RECT  116.545 0.52 116.805 5.815 ;
        RECT  117.13 190.585 117.33 191.315 ;
        RECT  118.075 0.17 118.845 0.43 ;
        RECT  118.075 0.17 118.335 11.5 ;
        RECT  118.585 0.17 118.845 11.5 ;
        RECT  117.625 190.585 117.825 191.315 ;
        RECT  118.125 190.585 118.325 191.315 ;
        RECT  118.625 190.585 118.825 191.315 ;
        RECT  120.115 0.17 120.885 0.43 ;
        RECT  120.115 0.17 120.375 10.48 ;
        RECT  120.625 0.17 120.885 10.99 ;
        RECT  119.12 190.585 119.32 191.315 ;
        RECT  119.94 190.585 120.14 191.315 ;
        RECT  121.135 0.17 121.905 0.94 ;
        RECT  121.135 0.17 121.395 8.7 ;
        RECT  121.645 0.17 121.905 12.9 ;
        RECT  120.435 190.585 120.635 191.315 ;
        RECT  120.935 190.585 121.135 191.315 ;
        RECT  121.435 190.585 121.635 191.315 ;
        RECT  121.93 190.585 122.13 191.315 ;
        RECT  122.155 0.52 122.415 2.485 ;
        RECT  122.75 190.585 122.95 191.315 ;
        RECT  123.02 0.52 123.28 14.11 ;
        RECT  123.245 190.585 123.445 191.315 ;
        RECT  123.53 0.52 123.79 2.335 ;
        RECT  123.745 190.585 123.945 191.315 ;
        RECT  124.245 190.585 124.445 191.315 ;
        RECT  124.74 190.585 124.94 191.315 ;
        RECT  126.93 0.52 127.19 5.16 ;
        RECT  126.41 4.9 127.19 5.16 ;
        RECT  126.41 4.9 126.67 6.64 ;
        RECT  125.56 190.585 125.76 191.315 ;
        RECT  126.055 190.585 126.255 191.315 ;
        RECT  126.555 190.585 126.755 191.315 ;
        RECT  127.055 190.585 127.255 191.315 ;
        RECT  127.55 190.585 127.75 191.315 ;
        RECT  128.295 0.17 129.065 0.94 ;
        RECT  128.295 0.17 128.555 12.9 ;
        RECT  128.805 0.17 129.065 12.9 ;
        RECT  127.785 0.52 128.045 5.815 ;
        RECT  128.37 190.585 128.57 191.315 ;
        RECT  129.315 0.17 130.085 0.43 ;
        RECT  129.315 0.17 129.575 11.5 ;
        RECT  129.825 0.17 130.085 11.5 ;
        RECT  128.865 190.585 129.065 191.315 ;
        RECT  129.365 190.585 129.565 191.315 ;
        RECT  129.865 190.585 130.065 191.315 ;
        RECT  131.355 0.17 132.125 0.43 ;
        RECT  131.355 0.17 131.615 10.48 ;
        RECT  131.865 0.17 132.125 10.99 ;
        RECT  130.36 190.585 130.56 191.315 ;
        RECT  131.18 190.585 131.38 191.315 ;
        RECT  132.375 0.17 133.145 0.94 ;
        RECT  132.375 0.17 132.635 8.7 ;
        RECT  132.885 0.17 133.145 12.9 ;
        RECT  131.675 190.585 131.875 191.315 ;
        RECT  132.175 190.585 132.375 191.315 ;
        RECT  132.675 190.585 132.875 191.315 ;
        RECT  133.17 190.585 133.37 191.315 ;
        RECT  133.395 0.52 133.655 2.485 ;
        RECT  133.99 190.585 134.19 191.315 ;
        RECT  134.26 0.52 134.52 14.11 ;
        RECT  134.485 190.585 134.685 191.315 ;
        RECT  134.77 0.52 135.03 2.335 ;
        RECT  134.985 190.585 135.185 191.315 ;
        RECT  135.485 190.585 135.685 191.315 ;
        RECT  135.98 190.585 136.18 191.315 ;
        RECT  138.17 0.52 138.43 5.16 ;
        RECT  137.65 4.9 138.43 5.16 ;
        RECT  137.65 4.9 137.91 6.64 ;
        RECT  136.8 190.585 137 191.315 ;
        RECT  137.295 190.585 137.495 191.315 ;
        RECT  137.795 190.585 137.995 191.315 ;
        RECT  138.295 190.585 138.495 191.315 ;
        RECT  138.79 190.585 138.99 191.315 ;
        RECT  139.535 0.17 140.305 0.94 ;
        RECT  139.535 0.17 139.795 12.9 ;
        RECT  140.045 0.17 140.305 12.9 ;
        RECT  139.025 0.52 139.285 5.815 ;
        RECT  139.61 190.585 139.81 191.315 ;
        RECT  140.555 0.17 141.325 0.43 ;
        RECT  140.555 0.17 140.815 11.5 ;
        RECT  141.065 0.17 141.325 11.5 ;
        RECT  140.105 190.585 140.305 191.315 ;
        RECT  140.605 190.585 140.805 191.315 ;
        RECT  141.105 190.585 141.305 191.315 ;
        RECT  142.595 0.17 143.365 0.43 ;
        RECT  142.595 0.17 142.855 10.48 ;
        RECT  143.105 0.17 143.365 10.99 ;
        RECT  141.6 190.585 141.8 191.315 ;
        RECT  142.42 190.585 142.62 191.315 ;
        RECT  143.615 0.17 144.385 0.94 ;
        RECT  143.615 0.17 143.875 8.7 ;
        RECT  144.125 0.17 144.385 12.9 ;
        RECT  142.915 190.585 143.115 191.315 ;
        RECT  143.415 190.585 143.615 191.315 ;
        RECT  143.915 190.585 144.115 191.315 ;
        RECT  144.41 190.585 144.61 191.315 ;
        RECT  144.635 0.52 144.895 2.485 ;
        RECT  145.23 190.585 145.43 191.315 ;
        RECT  145.5 0.52 145.76 14.11 ;
        RECT  145.725 190.585 145.925 191.315 ;
        RECT  146.01 0.52 146.27 2.335 ;
        RECT  146.225 190.585 146.425 191.315 ;
        RECT  146.725 190.585 146.925 191.315 ;
        RECT  147.22 190.585 147.42 191.315 ;
        RECT  149.41 0.52 149.67 5.16 ;
        RECT  148.89 4.9 149.67 5.16 ;
        RECT  148.89 4.9 149.15 6.64 ;
        RECT  148.04 190.585 148.24 191.315 ;
        RECT  148.535 190.585 148.735 191.315 ;
        RECT  149.035 190.585 149.235 191.315 ;
        RECT  149.535 190.585 149.735 191.315 ;
        RECT  150.03 190.585 150.23 191.315 ;
        RECT  150.775 0.17 151.545 0.94 ;
        RECT  150.775 0.17 151.035 12.9 ;
        RECT  151.285 0.17 151.545 12.9 ;
        RECT  150.265 0.52 150.525 5.815 ;
        RECT  150.85 190.585 151.05 191.315 ;
        RECT  151.795 0.17 152.565 0.43 ;
        RECT  151.795 0.17 152.055 11.5 ;
        RECT  152.305 0.17 152.565 11.5 ;
        RECT  151.345 190.585 151.545 191.315 ;
        RECT  151.845 190.585 152.045 191.315 ;
        RECT  152.345 190.585 152.545 191.315 ;
        RECT  153.835 0.17 154.605 0.43 ;
        RECT  153.835 0.17 154.095 10.48 ;
        RECT  154.345 0.17 154.605 10.99 ;
        RECT  152.84 190.585 153.04 191.315 ;
        RECT  153.66 190.585 153.86 191.315 ;
        RECT  154.855 0.17 155.625 0.94 ;
        RECT  154.855 0.17 155.115 8.7 ;
        RECT  155.365 0.17 155.625 12.9 ;
        RECT  154.155 190.585 154.355 191.315 ;
        RECT  154.655 190.585 154.855 191.315 ;
        RECT  155.155 190.585 155.355 191.315 ;
        RECT  155.65 190.585 155.85 191.315 ;
        RECT  155.875 0.52 156.135 2.485 ;
        RECT  156.47 190.585 156.67 191.315 ;
        RECT  156.74 0.52 157 14.11 ;
        RECT  156.965 190.585 157.165 191.315 ;
        RECT  157.25 0.52 157.51 2.335 ;
        RECT  157.465 190.585 157.665 191.315 ;
        RECT  157.965 190.585 158.165 191.315 ;
        RECT  158.46 190.585 158.66 191.315 ;
        RECT  160.65 0.52 160.91 5.16 ;
        RECT  160.13 4.9 160.91 5.16 ;
        RECT  160.13 4.9 160.39 6.64 ;
        RECT  159.28 190.585 159.48 191.315 ;
        RECT  159.775 190.585 159.975 191.315 ;
        RECT  160.275 190.585 160.475 191.315 ;
        RECT  160.775 190.585 160.975 191.315 ;
        RECT  161.27 190.585 161.47 191.315 ;
        RECT  162.015 0.17 162.785 0.94 ;
        RECT  162.015 0.17 162.275 12.9 ;
        RECT  162.525 0.17 162.785 12.9 ;
        RECT  161.505 0.52 161.765 5.815 ;
        RECT  162.09 190.585 162.29 191.315 ;
        RECT  163.035 0.17 163.805 0.43 ;
        RECT  163.035 0.17 163.295 11.5 ;
        RECT  163.545 0.17 163.805 11.5 ;
        RECT  162.585 190.585 162.785 191.315 ;
        RECT  163.085 190.585 163.285 191.315 ;
        RECT  163.585 190.585 163.785 191.315 ;
        RECT  165.075 0.17 165.845 0.43 ;
        RECT  165.075 0.17 165.335 10.48 ;
        RECT  165.585 0.17 165.845 10.99 ;
        RECT  164.08 190.585 164.28 191.315 ;
        RECT  164.9 190.585 165.1 191.315 ;
        RECT  166.095 0.17 166.865 0.94 ;
        RECT  166.095 0.17 166.355 8.7 ;
        RECT  166.605 0.17 166.865 12.9 ;
        RECT  165.395 190.585 165.595 191.315 ;
        RECT  165.895 190.585 166.095 191.315 ;
        RECT  166.395 190.585 166.595 191.315 ;
        RECT  166.89 190.585 167.09 191.315 ;
        RECT  167.115 0.52 167.375 2.485 ;
        RECT  167.71 190.585 167.91 191.315 ;
        RECT  167.98 0.52 168.24 14.11 ;
        RECT  168.205 190.585 168.405 191.315 ;
        RECT  168.49 0.52 168.75 2.335 ;
        RECT  168.705 190.585 168.905 191.315 ;
        RECT  169.205 190.585 169.405 191.315 ;
        RECT  169.7 190.585 169.9 191.315 ;
        RECT  171.89 0.52 172.15 5.16 ;
        RECT  171.37 4.9 172.15 5.16 ;
        RECT  171.37 4.9 171.63 6.64 ;
        RECT  170.52 190.585 170.72 191.315 ;
        RECT  171.015 190.585 171.215 191.315 ;
        RECT  171.515 190.585 171.715 191.315 ;
        RECT  172.015 190.585 172.215 191.315 ;
        RECT  172.51 190.585 172.71 191.315 ;
        RECT  173.255 0.17 174.025 0.94 ;
        RECT  173.255 0.17 173.515 12.9 ;
        RECT  173.765 0.17 174.025 12.9 ;
        RECT  172.745 0.52 173.005 5.815 ;
        RECT  173.33 190.585 173.53 191.315 ;
        RECT  174.275 0.17 175.045 0.43 ;
        RECT  174.275 0.17 174.535 11.5 ;
        RECT  174.785 0.17 175.045 11.5 ;
        RECT  173.825 190.585 174.025 191.315 ;
        RECT  174.325 190.585 174.525 191.315 ;
        RECT  174.825 190.585 175.025 191.315 ;
        RECT  176.315 0.17 177.085 0.43 ;
        RECT  176.315 0.17 176.575 10.48 ;
        RECT  176.825 0.17 177.085 10.99 ;
        RECT  175.32 190.585 175.52 191.315 ;
        RECT  176.14 190.585 176.34 191.315 ;
        RECT  177.335 0.17 178.105 0.94 ;
        RECT  177.335 0.17 177.595 8.7 ;
        RECT  177.845 0.17 178.105 12.9 ;
        RECT  176.635 190.585 176.835 191.315 ;
        RECT  177.135 190.585 177.335 191.315 ;
        RECT  177.635 190.585 177.835 191.315 ;
        RECT  178.13 190.585 178.33 191.315 ;
        RECT  178.355 0.52 178.615 2.485 ;
        RECT  178.95 190.585 179.15 191.315 ;
        RECT  179.22 0.52 179.48 14.11 ;
        RECT  179.445 190.585 179.645 191.315 ;
        RECT  179.73 0.52 179.99 2.335 ;
        RECT  179.945 190.585 180.145 191.315 ;
        RECT  180.445 190.585 180.645 191.315 ;
        RECT  182.435 0.17 183.205 0.43 ;
        RECT  182.435 0.17 182.695 8.7 ;
        RECT  182.945 0.17 183.205 8.7 ;
        RECT  183.455 0.17 184.225 0.94 ;
        RECT  183.455 0.17 183.715 8.7 ;
        RECT  183.965 0.17 184.225 8.7 ;
        RECT  184.475 0.17 185.245 0.43 ;
        RECT  184.475 0.17 184.735 8.7 ;
        RECT  184.985 0.17 185.245 8.7 ;
        RECT  185.495 0.17 186.265 0.94 ;
        RECT  185.495 0.17 185.755 8.7 ;
        RECT  186.005 0.17 186.265 8.7 ;
        RECT  186.515 0.17 187.285 0.43 ;
        RECT  186.515 0.17 186.775 8.7 ;
        RECT  187.025 0.17 187.285 8.7 ;
        RECT  187.535 0.17 188.305 0.94 ;
        RECT  187.535 0.17 187.795 8.7 ;
        RECT  188.045 0.17 188.305 8.7 ;
        RECT  180.94 190.585 181.14 191.315 ;
        RECT  181.76 190.585 181.96 191.315 ;
        RECT  182.755 190.585 182.955 191.315 ;
        RECT  190.24 0.17 191.01 0.94 ;
        RECT  190.24 0.17 190.5 8.7 ;
        RECT  190.75 0.17 191.01 8.7 ;
        RECT  188.71 0.3 188.97 8.7 ;
        RECT  189.22 0 189.48 8.7 ;
        RECT  189.73 0 189.99 8.7 ;
        RECT  191.26 0 191.52 8.7 ;
        RECT  191.77 0 192.03 8.7 ;
        RECT  192.28 0.52 192.54 8.7 ;
        RECT  192.79 0.52 193.05 8.7 ;
        RECT  193.3 0.52 193.56 8.7 ;
        RECT  195.34 0.17 196.11 0.94 ;
        RECT  195.34 0.17 195.6 8.7 ;
        RECT  195.85 0.17 196.11 8.7 ;
        RECT  196.36 0.17 197.13 0.43 ;
        RECT  196.36 0.17 196.62 8.7 ;
        RECT  196.87 0.17 197.13 8.7 ;
        RECT  193.81 0.52 194.07 8.7 ;
        RECT  194.32 0 194.58 8.7 ;
        RECT  194.83 0 195.09 8.7 ;
        RECT  197.38 0.3 197.64 8.7 ;
        RECT  197.89 0.3 198.15 8.7 ;
        RECT  199.93 0.17 200.7 0.94 ;
        RECT  199.93 0.17 200.19 8.7 ;
        RECT  200.44 0.17 200.7 8.7 ;
        RECT  198.4 0.3 198.66 8.7 ;
        RECT  198.91 0.3 199.17 8.7 ;
        RECT  199.42 0.3 199.68 8.7 ;
        RECT  200.95 0.52 201.21 8.7 ;
        RECT  201.46 0.52 201.72 8.7 ;
        RECT  201.97 0.3 202.23 8.7 ;
        RECT  202.48 0.52 202.74 8.7 ;
        RECT  202.99 0.52 203.25 8.7 ;
        RECT  203.5 0.3 203.76 8.7 ;
        RECT  204.01 0.52 204.27 8.7 ;
        RECT  204.52 0.52 204.78 8.7 ;
        RECT  205.03 0.52 205.29 8.7 ;
        RECT  205.54 0.52 205.8 8.7 ;
        RECT  206.05 0.52 206.31 8.7 ;
        RECT  206.56 0.3 206.82 8.7 ;
        RECT  207.07 0.52 207.33 8.7 ;
        RECT  207.58 0.52 207.84 8.7 ;
        RECT  208.09 0.3 208.35 8.7 ;
        RECT  210.13 0.17 210.9 0.94 ;
        RECT  210.13 0.17 210.39 8.7 ;
        RECT  210.64 0.17 210.9 8.7 ;
        RECT  208.6 0.52 208.86 8.7 ;
        RECT  209.11 0.52 209.37 8.7 ;
        RECT  209.62 0.3 209.88 8.7 ;
        RECT  211.15 0.52 211.41 8.7 ;
        RECT  211.66 0.52 211.92 8.7 ;
        RECT  212.17 0.52 212.43 8.7 ;
        RECT  212.68 0.52 212.94 8.7 ;
        RECT  213.19 0.52 213.45 8.7 ;
        RECT  213.7 0.52 213.96 8.7 ;
        RECT  214.21 0.52 214.47 8.7 ;
        RECT  216.25 0.17 217.02 0.94 ;
        RECT  216.25 0.17 216.51 8.7 ;
        RECT  216.76 0.17 217.02 8.7 ;
        RECT  214.72 0.52 214.98 8.7 ;
        RECT  215.23 0 215.49 8.7 ;
        RECT  215.74 0 216 8.7 ;
        RECT  217.27 0 217.53 8.7 ;
        RECT  219.31 0.17 220.08 0.43 ;
        RECT  219.31 0.17 219.57 8.7 ;
        RECT  219.82 0.17 220.08 8.7 ;
        RECT  217.78 0 218.04 8.7 ;
        RECT  218.29 0.3 218.55 8.7 ;
        RECT  218.8 0.3 219.06 8.7 ;
        RECT  220.33 0.3 220.59 8.7 ;
        RECT  220.84 0.3 221.1 8.7 ;
        RECT  221.35 0.3 221.61 8.7 ;
        RECT  221.86 0.3 222.12 8.7 ;
        RECT  222.37 0.52 222.63 8.7 ;
        RECT  222.88 0.52 223.14 8.7 ;
        RECT  224.92 0.17 225.69 0.43 ;
        RECT  224.92 0.17 225.18 8.7 ;
        RECT  225.43 0.17 225.69 8.7 ;
        RECT  225.94 0.17 226.71 0.94 ;
        RECT  225.94 0.17 226.2 25.5 ;
        RECT  226.45 0.17 226.71 33.9 ;
        RECT  226.96 0.17 227.73 0.43 ;
        RECT  226.96 0.17 227.22 8.7 ;
        RECT  227.47 0.17 227.73 8.7 ;
        RECT  228.335 0.17 229.105 0.94 ;
        RECT  228.335 0.17 228.595 8.7 ;
        RECT  228.845 0.17 229.105 8.7 ;
        RECT  229.355 0.17 230.125 0.43 ;
        RECT  229.355 0.17 229.615 8.7 ;
        RECT  229.865 0.17 230.125 8.7 ;
        RECT  230.375 0.17 231.145 0.94 ;
        RECT  230.375 0.17 230.635 8.7 ;
        RECT  230.885 0.17 231.145 8.7 ;
        RECT  231.395 0.17 232.165 0.43 ;
        RECT  231.395 0.17 231.655 8.7 ;
        RECT  231.905 0.17 232.165 8.7 ;
        RECT  232.415 0.17 233.185 0.94 ;
        RECT  232.415 0.17 232.675 8.7 ;
        RECT  232.925 0.17 233.185 8.7 ;
        RECT  223.39 0.3 223.65 8.7 ;
        RECT  233.435 0.17 234.205 0.43 ;
        RECT  233.435 0.17 233.695 8.7 ;
        RECT  233.945 0.17 234.205 8.7 ;
        RECT  223.9 0.3 224.16 8.7 ;
        RECT  224.41 0.52 224.67 8.7 ;
        RECT  233.685 190.585 233.885 191.315 ;
        RECT  234.68 190.585 234.88 191.315 ;
        RECT  235.5 190.585 235.7 191.315 ;
        RECT  235.995 190.585 236.195 191.315 ;
        RECT  236.495 190.585 236.695 191.315 ;
        RECT  236.65 0.52 236.91 2.335 ;
        RECT  236.995 190.585 237.195 191.315 ;
        RECT  237.16 0.52 237.42 14.11 ;
        RECT  237.49 190.585 237.69 191.315 ;
        RECT  238.535 0.17 239.305 0.94 ;
        RECT  239.045 0.17 239.305 8.7 ;
        RECT  238.535 0.17 238.795 12.9 ;
        RECT  238.025 0.52 238.285 2.485 ;
        RECT  238.31 190.585 238.51 191.315 ;
        RECT  239.555 0.17 240.325 0.43 ;
        RECT  240.065 0.17 240.325 10.48 ;
        RECT  239.555 0.17 239.815 10.99 ;
        RECT  238.805 190.585 239.005 191.315 ;
        RECT  239.305 190.585 239.505 191.315 ;
        RECT  239.805 190.585 240.005 191.315 ;
        RECT  240.3 190.585 240.5 191.315 ;
        RECT  241.595 0.17 242.365 0.43 ;
        RECT  241.595 0.17 241.855 11.5 ;
        RECT  242.105 0.17 242.365 11.5 ;
        RECT  241.12 190.585 241.32 191.315 ;
        RECT  241.615 190.585 241.815 191.315 ;
        RECT  242.615 0.17 243.385 0.94 ;
        RECT  242.615 0.17 242.875 12.9 ;
        RECT  243.125 0.17 243.385 12.9 ;
        RECT  242.115 190.585 242.315 191.315 ;
        RECT  242.615 190.585 242.815 191.315 ;
        RECT  243.11 190.585 243.31 191.315 ;
        RECT  243.635 0.52 243.895 5.815 ;
        RECT  244.49 0.52 244.75 5.16 ;
        RECT  244.49 4.9 245.27 5.16 ;
        RECT  245.01 4.9 245.27 6.64 ;
        RECT  243.93 190.585 244.13 191.315 ;
        RECT  244.425 190.585 244.625 191.315 ;
        RECT  244.925 190.585 245.125 191.315 ;
        RECT  245.425 190.585 245.625 191.315 ;
        RECT  245.92 190.585 246.12 191.315 ;
        RECT  246.74 190.585 246.94 191.315 ;
        RECT  247.235 190.585 247.435 191.315 ;
        RECT  247.735 190.585 247.935 191.315 ;
        RECT  247.89 0.52 248.15 2.335 ;
        RECT  248.235 190.585 248.435 191.315 ;
        RECT  248.4 0.52 248.66 14.11 ;
        RECT  248.73 190.585 248.93 191.315 ;
        RECT  249.775 0.17 250.545 0.94 ;
        RECT  250.285 0.17 250.545 8.7 ;
        RECT  249.775 0.17 250.035 12.9 ;
        RECT  249.265 0.52 249.525 2.485 ;
        RECT  249.55 190.585 249.75 191.315 ;
        RECT  250.795 0.17 251.565 0.43 ;
        RECT  251.305 0.17 251.565 10.48 ;
        RECT  250.795 0.17 251.055 10.99 ;
        RECT  250.045 190.585 250.245 191.315 ;
        RECT  250.545 190.585 250.745 191.315 ;
        RECT  251.045 190.585 251.245 191.315 ;
        RECT  251.54 190.585 251.74 191.315 ;
        RECT  252.835 0.17 253.605 0.43 ;
        RECT  252.835 0.17 253.095 11.5 ;
        RECT  253.345 0.17 253.605 11.5 ;
        RECT  252.36 190.585 252.56 191.315 ;
        RECT  252.855 190.585 253.055 191.315 ;
        RECT  253.855 0.17 254.625 0.94 ;
        RECT  253.855 0.17 254.115 12.9 ;
        RECT  254.365 0.17 254.625 12.9 ;
        RECT  253.355 190.585 253.555 191.315 ;
        RECT  253.855 190.585 254.055 191.315 ;
        RECT  254.35 190.585 254.55 191.315 ;
        RECT  254.875 0.52 255.135 5.815 ;
        RECT  255.73 0.52 255.99 5.16 ;
        RECT  255.73 4.9 256.51 5.16 ;
        RECT  256.25 4.9 256.51 6.64 ;
        RECT  255.17 190.585 255.37 191.315 ;
        RECT  255.665 190.585 255.865 191.315 ;
        RECT  256.165 190.585 256.365 191.315 ;
        RECT  256.665 190.585 256.865 191.315 ;
        RECT  257.16 190.585 257.36 191.315 ;
        RECT  257.98 190.585 258.18 191.315 ;
        RECT  258.475 190.585 258.675 191.315 ;
        RECT  258.975 190.585 259.175 191.315 ;
        RECT  259.13 0.52 259.39 2.335 ;
        RECT  259.475 190.585 259.675 191.315 ;
        RECT  259.64 0.52 259.9 14.11 ;
        RECT  259.97 190.585 260.17 191.315 ;
        RECT  261.015 0.17 261.785 0.94 ;
        RECT  261.525 0.17 261.785 8.7 ;
        RECT  261.015 0.17 261.275 12.9 ;
        RECT  260.505 0.52 260.765 2.485 ;
        RECT  260.79 190.585 260.99 191.315 ;
        RECT  262.035 0.17 262.805 0.43 ;
        RECT  262.545 0.17 262.805 10.48 ;
        RECT  262.035 0.17 262.295 10.99 ;
        RECT  261.285 190.585 261.485 191.315 ;
        RECT  261.785 190.585 261.985 191.315 ;
        RECT  262.285 190.585 262.485 191.315 ;
        RECT  262.78 190.585 262.98 191.315 ;
        RECT  264.075 0.17 264.845 0.43 ;
        RECT  264.075 0.17 264.335 11.5 ;
        RECT  264.585 0.17 264.845 11.5 ;
        RECT  263.6 190.585 263.8 191.315 ;
        RECT  264.095 190.585 264.295 191.315 ;
        RECT  265.095 0.17 265.865 0.94 ;
        RECT  265.095 0.17 265.355 12.9 ;
        RECT  265.605 0.17 265.865 12.9 ;
        RECT  264.595 190.585 264.795 191.315 ;
        RECT  265.095 190.585 265.295 191.315 ;
        RECT  265.59 190.585 265.79 191.315 ;
        RECT  266.115 0.52 266.375 5.815 ;
        RECT  266.97 0.52 267.23 5.16 ;
        RECT  266.97 4.9 267.75 5.16 ;
        RECT  267.49 4.9 267.75 6.64 ;
        RECT  266.41 190.585 266.61 191.315 ;
        RECT  266.905 190.585 267.105 191.315 ;
        RECT  267.405 190.585 267.605 191.315 ;
        RECT  267.905 190.585 268.105 191.315 ;
        RECT  268.4 190.585 268.6 191.315 ;
        RECT  269.22 190.585 269.42 191.315 ;
        RECT  269.715 190.585 269.915 191.315 ;
        RECT  270.215 190.585 270.415 191.315 ;
        RECT  270.37 0.52 270.63 2.335 ;
        RECT  270.715 190.585 270.915 191.315 ;
        RECT  270.88 0.52 271.14 14.11 ;
        RECT  271.21 190.585 271.41 191.315 ;
        RECT  272.255 0.17 273.025 0.94 ;
        RECT  272.765 0.17 273.025 8.7 ;
        RECT  272.255 0.17 272.515 12.9 ;
        RECT  271.745 0.52 272.005 2.485 ;
        RECT  272.03 190.585 272.23 191.315 ;
        RECT  273.275 0.17 274.045 0.43 ;
        RECT  273.785 0.17 274.045 10.48 ;
        RECT  273.275 0.17 273.535 10.99 ;
        RECT  272.525 190.585 272.725 191.315 ;
        RECT  273.025 190.585 273.225 191.315 ;
        RECT  273.525 190.585 273.725 191.315 ;
        RECT  274.02 190.585 274.22 191.315 ;
        RECT  275.315 0.17 276.085 0.43 ;
        RECT  275.315 0.17 275.575 11.5 ;
        RECT  275.825 0.17 276.085 11.5 ;
        RECT  274.84 190.585 275.04 191.315 ;
        RECT  275.335 190.585 275.535 191.315 ;
        RECT  276.335 0.17 277.105 0.94 ;
        RECT  276.335 0.17 276.595 12.9 ;
        RECT  276.845 0.17 277.105 12.9 ;
        RECT  275.835 190.585 276.035 191.315 ;
        RECT  276.335 190.585 276.535 191.315 ;
        RECT  276.83 190.585 277.03 191.315 ;
        RECT  277.355 0.52 277.615 5.815 ;
        RECT  278.21 0.52 278.47 5.16 ;
        RECT  278.21 4.9 278.99 5.16 ;
        RECT  278.73 4.9 278.99 6.64 ;
        RECT  277.65 190.585 277.85 191.315 ;
        RECT  278.145 190.585 278.345 191.315 ;
        RECT  278.645 190.585 278.845 191.315 ;
        RECT  279.145 190.585 279.345 191.315 ;
        RECT  279.64 190.585 279.84 191.315 ;
        RECT  280.46 190.585 280.66 191.315 ;
        RECT  280.955 190.585 281.155 191.315 ;
        RECT  281.455 190.585 281.655 191.315 ;
        RECT  281.61 0.52 281.87 2.335 ;
        RECT  281.955 190.585 282.155 191.315 ;
        RECT  282.12 0.52 282.38 14.11 ;
        RECT  282.45 190.585 282.65 191.315 ;
        RECT  283.495 0.17 284.265 0.94 ;
        RECT  284.005 0.17 284.265 8.7 ;
        RECT  283.495 0.17 283.755 12.9 ;
        RECT  282.985 0.52 283.245 2.485 ;
        RECT  283.27 190.585 283.47 191.315 ;
        RECT  284.515 0.17 285.285 0.43 ;
        RECT  285.025 0.17 285.285 10.48 ;
        RECT  284.515 0.17 284.775 10.99 ;
        RECT  283.765 190.585 283.965 191.315 ;
        RECT  284.265 190.585 284.465 191.315 ;
        RECT  284.765 190.585 284.965 191.315 ;
        RECT  285.26 190.585 285.46 191.315 ;
        RECT  286.555 0.17 287.325 0.43 ;
        RECT  286.555 0.17 286.815 11.5 ;
        RECT  287.065 0.17 287.325 11.5 ;
        RECT  286.08 190.585 286.28 191.315 ;
        RECT  286.575 190.585 286.775 191.315 ;
        RECT  287.575 0.17 288.345 0.94 ;
        RECT  287.575 0.17 287.835 12.9 ;
        RECT  288.085 0.17 288.345 12.9 ;
        RECT  287.075 190.585 287.275 191.315 ;
        RECT  287.575 190.585 287.775 191.315 ;
        RECT  288.07 190.585 288.27 191.315 ;
        RECT  288.595 0.52 288.855 5.815 ;
        RECT  289.45 0.52 289.71 5.16 ;
        RECT  289.45 4.9 290.23 5.16 ;
        RECT  289.97 4.9 290.23 6.64 ;
        RECT  288.89 190.585 289.09 191.315 ;
        RECT  289.385 190.585 289.585 191.315 ;
        RECT  289.885 190.585 290.085 191.315 ;
        RECT  290.385 190.585 290.585 191.315 ;
        RECT  290.88 190.585 291.08 191.315 ;
        RECT  291.7 190.585 291.9 191.315 ;
        RECT  292.195 190.585 292.395 191.315 ;
        RECT  292.695 190.585 292.895 191.315 ;
        RECT  292.85 0.52 293.11 2.335 ;
        RECT  293.195 190.585 293.395 191.315 ;
        RECT  293.36 0.52 293.62 14.11 ;
        RECT  293.69 190.585 293.89 191.315 ;
        RECT  294.735 0.17 295.505 0.94 ;
        RECT  295.245 0.17 295.505 8.7 ;
        RECT  294.735 0.17 294.995 12.9 ;
        RECT  294.225 0.52 294.485 2.485 ;
        RECT  294.51 190.585 294.71 191.315 ;
        RECT  295.755 0.17 296.525 0.43 ;
        RECT  296.265 0.17 296.525 10.48 ;
        RECT  295.755 0.17 296.015 10.99 ;
        RECT  295.005 190.585 295.205 191.315 ;
        RECT  295.505 190.585 295.705 191.315 ;
        RECT  296.005 190.585 296.205 191.315 ;
        RECT  296.5 190.585 296.7 191.315 ;
        RECT  297.795 0.17 298.565 0.43 ;
        RECT  297.795 0.17 298.055 11.5 ;
        RECT  298.305 0.17 298.565 11.5 ;
        RECT  297.32 190.585 297.52 191.315 ;
        RECT  297.815 190.585 298.015 191.315 ;
        RECT  298.815 0.17 299.585 0.94 ;
        RECT  298.815 0.17 299.075 12.9 ;
        RECT  299.325 0.17 299.585 12.9 ;
        RECT  298.315 190.585 298.515 191.315 ;
        RECT  298.815 190.585 299.015 191.315 ;
        RECT  299.31 190.585 299.51 191.315 ;
        RECT  299.835 0.52 300.095 5.815 ;
        RECT  300.69 0.52 300.95 5.16 ;
        RECT  300.69 4.9 301.47 5.16 ;
        RECT  301.21 4.9 301.47 6.64 ;
        RECT  300.13 190.585 300.33 191.315 ;
        RECT  300.625 190.585 300.825 191.315 ;
        RECT  301.125 190.585 301.325 191.315 ;
        RECT  301.625 190.585 301.825 191.315 ;
        RECT  302.12 190.585 302.32 191.315 ;
        RECT  302.94 190.585 303.14 191.315 ;
        RECT  303.435 190.585 303.635 191.315 ;
        RECT  303.935 190.585 304.135 191.315 ;
        RECT  304.09 0.52 304.35 2.335 ;
        RECT  304.435 190.585 304.635 191.315 ;
        RECT  304.6 0.52 304.86 14.11 ;
        RECT  304.93 190.585 305.13 191.315 ;
        RECT  305.975 0.17 306.745 0.94 ;
        RECT  306.485 0.17 306.745 8.7 ;
        RECT  305.975 0.17 306.235 12.9 ;
        RECT  305.465 0.52 305.725 2.485 ;
        RECT  305.75 190.585 305.95 191.315 ;
        RECT  306.995 0.17 307.765 0.43 ;
        RECT  307.505 0.17 307.765 10.48 ;
        RECT  306.995 0.17 307.255 10.99 ;
        RECT  306.245 190.585 306.445 191.315 ;
        RECT  306.745 190.585 306.945 191.315 ;
        RECT  307.245 190.585 307.445 191.315 ;
        RECT  307.74 190.585 307.94 191.315 ;
        RECT  309.035 0.17 309.805 0.43 ;
        RECT  309.035 0.17 309.295 11.5 ;
        RECT  309.545 0.17 309.805 11.5 ;
        RECT  308.56 190.585 308.76 191.315 ;
        RECT  309.055 190.585 309.255 191.315 ;
        RECT  310.055 0.17 310.825 0.94 ;
        RECT  310.055 0.17 310.315 12.9 ;
        RECT  310.565 0.17 310.825 12.9 ;
        RECT  309.555 190.585 309.755 191.315 ;
        RECT  310.055 190.585 310.255 191.315 ;
        RECT  310.55 190.585 310.75 191.315 ;
        RECT  311.075 0.52 311.335 5.815 ;
        RECT  311.93 0.52 312.19 5.16 ;
        RECT  311.93 4.9 312.71 5.16 ;
        RECT  312.45 4.9 312.71 6.64 ;
        RECT  311.37 190.585 311.57 191.315 ;
        RECT  311.865 190.585 312.065 191.315 ;
        RECT  312.365 190.585 312.565 191.315 ;
        RECT  312.865 190.585 313.065 191.315 ;
        RECT  313.36 190.585 313.56 191.315 ;
        RECT  314.18 190.585 314.38 191.315 ;
        RECT  314.675 190.585 314.875 191.315 ;
        RECT  315.175 190.585 315.375 191.315 ;
        RECT  315.33 0.52 315.59 2.335 ;
        RECT  315.675 190.585 315.875 191.315 ;
        RECT  315.84 0.52 316.1 14.11 ;
        RECT  316.17 190.585 316.37 191.315 ;
        RECT  317.215 0.17 317.985 0.94 ;
        RECT  317.725 0.17 317.985 8.7 ;
        RECT  317.215 0.17 317.475 12.9 ;
        RECT  316.705 0.52 316.965 2.485 ;
        RECT  316.99 190.585 317.19 191.315 ;
        RECT  318.235 0.17 319.005 0.43 ;
        RECT  318.745 0.17 319.005 10.48 ;
        RECT  318.235 0.17 318.495 10.99 ;
        RECT  317.485 190.585 317.685 191.315 ;
        RECT  317.985 190.585 318.185 191.315 ;
        RECT  318.485 190.585 318.685 191.315 ;
        RECT  318.98 190.585 319.18 191.315 ;
        RECT  320.275 0.17 321.045 0.43 ;
        RECT  320.275 0.17 320.535 11.5 ;
        RECT  320.785 0.17 321.045 11.5 ;
        RECT  319.8 190.585 320 191.315 ;
        RECT  320.295 190.585 320.495 191.315 ;
        RECT  321.295 0.17 322.065 0.94 ;
        RECT  321.295 0.17 321.555 12.9 ;
        RECT  321.805 0.17 322.065 12.9 ;
        RECT  320.795 190.585 320.995 191.315 ;
        RECT  321.295 190.585 321.495 191.315 ;
        RECT  321.79 190.585 321.99 191.315 ;
        RECT  322.315 0.52 322.575 5.815 ;
        RECT  323.17 0.52 323.43 5.16 ;
        RECT  323.17 4.9 323.95 5.16 ;
        RECT  323.69 4.9 323.95 6.64 ;
        RECT  322.61 190.585 322.81 191.315 ;
        RECT  323.105 190.585 323.305 191.315 ;
        RECT  323.605 190.585 323.805 191.315 ;
        RECT  324.105 190.585 324.305 191.315 ;
        RECT  324.6 190.585 324.8 191.315 ;
        RECT  325.42 190.585 325.62 191.315 ;
        RECT  325.915 190.585 326.115 191.315 ;
        RECT  326.415 190.585 326.615 191.315 ;
        RECT  326.57 0.52 326.83 2.335 ;
        RECT  326.915 190.585 327.115 191.315 ;
        RECT  327.08 0.52 327.34 14.11 ;
        RECT  327.41 190.585 327.61 191.315 ;
        RECT  328.455 0.17 329.225 0.94 ;
        RECT  328.965 0.17 329.225 8.7 ;
        RECT  328.455 0.17 328.715 12.9 ;
        RECT  327.945 0.52 328.205 2.485 ;
        RECT  328.23 190.585 328.43 191.315 ;
        RECT  329.475 0.17 330.245 0.43 ;
        RECT  329.985 0.17 330.245 10.48 ;
        RECT  329.475 0.17 329.735 10.99 ;
        RECT  328.725 190.585 328.925 191.315 ;
        RECT  329.225 190.585 329.425 191.315 ;
        RECT  329.725 190.585 329.925 191.315 ;
        RECT  330.22 190.585 330.42 191.315 ;
        RECT  331.515 0.17 332.285 0.43 ;
        RECT  331.515 0.17 331.775 11.5 ;
        RECT  332.025 0.17 332.285 11.5 ;
        RECT  331.04 190.585 331.24 191.315 ;
        RECT  331.535 190.585 331.735 191.315 ;
        RECT  332.535 0.17 333.305 0.94 ;
        RECT  332.535 0.17 332.795 12.9 ;
        RECT  333.045 0.17 333.305 12.9 ;
        RECT  332.035 190.585 332.235 191.315 ;
        RECT  332.535 190.585 332.735 191.315 ;
        RECT  333.03 190.585 333.23 191.315 ;
        RECT  333.555 0.52 333.815 5.815 ;
        RECT  334.41 0.52 334.67 5.16 ;
        RECT  334.41 4.9 335.19 5.16 ;
        RECT  334.93 4.9 335.19 6.64 ;
        RECT  333.85 190.585 334.05 191.315 ;
        RECT  334.345 190.585 334.545 191.315 ;
        RECT  334.845 190.585 335.045 191.315 ;
        RECT  335.345 190.585 335.545 191.315 ;
        RECT  335.84 190.585 336.04 191.315 ;
        RECT  336.66 190.585 336.86 191.315 ;
        RECT  337.155 190.585 337.355 191.315 ;
        RECT  337.655 190.585 337.855 191.315 ;
        RECT  337.81 0.52 338.07 2.335 ;
        RECT  338.155 190.585 338.355 191.315 ;
        RECT  338.32 0.52 338.58 14.11 ;
        RECT  338.65 190.585 338.85 191.315 ;
        RECT  339.695 0.17 340.465 0.94 ;
        RECT  340.205 0.17 340.465 8.7 ;
        RECT  339.695 0.17 339.955 12.9 ;
        RECT  339.185 0.52 339.445 2.485 ;
        RECT  339.47 190.585 339.67 191.315 ;
        RECT  340.715 0.17 341.485 0.43 ;
        RECT  341.225 0.17 341.485 10.48 ;
        RECT  340.715 0.17 340.975 10.99 ;
        RECT  339.965 190.585 340.165 191.315 ;
        RECT  340.465 190.585 340.665 191.315 ;
        RECT  340.965 190.585 341.165 191.315 ;
        RECT  341.46 190.585 341.66 191.315 ;
        RECT  342.755 0.17 343.525 0.43 ;
        RECT  342.755 0.17 343.015 11.5 ;
        RECT  343.265 0.17 343.525 11.5 ;
        RECT  342.28 190.585 342.48 191.315 ;
        RECT  342.775 190.585 342.975 191.315 ;
        RECT  343.775 0.17 344.545 0.94 ;
        RECT  343.775 0.17 344.035 12.9 ;
        RECT  344.285 0.17 344.545 12.9 ;
        RECT  343.275 190.585 343.475 191.315 ;
        RECT  343.775 190.585 343.975 191.315 ;
        RECT  344.27 190.585 344.47 191.315 ;
        RECT  344.795 0.52 345.055 5.815 ;
        RECT  345.65 0.52 345.91 5.16 ;
        RECT  345.65 4.9 346.43 5.16 ;
        RECT  346.17 4.9 346.43 6.64 ;
        RECT  345.09 190.585 345.29 191.315 ;
        RECT  345.585 190.585 345.785 191.315 ;
        RECT  346.085 190.585 346.285 191.315 ;
        RECT  346.585 190.585 346.785 191.315 ;
        RECT  347.08 190.585 347.28 191.315 ;
        RECT  347.9 190.585 348.1 191.315 ;
        RECT  348.395 190.585 348.595 191.315 ;
        RECT  348.895 190.585 349.095 191.315 ;
        RECT  349.05 0.52 349.31 2.335 ;
        RECT  349.395 190.585 349.595 191.315 ;
        RECT  349.56 0.52 349.82 14.11 ;
        RECT  349.89 190.585 350.09 191.315 ;
        RECT  350.935 0.17 351.705 0.94 ;
        RECT  351.445 0.17 351.705 8.7 ;
        RECT  350.935 0.17 351.195 12.9 ;
        RECT  350.425 0.52 350.685 2.485 ;
        RECT  350.71 190.585 350.91 191.315 ;
        RECT  351.955 0.17 352.725 0.43 ;
        RECT  352.465 0.17 352.725 10.48 ;
        RECT  351.955 0.17 352.215 10.99 ;
        RECT  351.205 190.585 351.405 191.315 ;
        RECT  351.705 190.585 351.905 191.315 ;
        RECT  352.205 190.585 352.405 191.315 ;
        RECT  352.7 190.585 352.9 191.315 ;
        RECT  353.995 0.17 354.765 0.43 ;
        RECT  353.995 0.17 354.255 11.5 ;
        RECT  354.505 0.17 354.765 11.5 ;
        RECT  353.52 190.585 353.72 191.315 ;
        RECT  354.015 190.585 354.215 191.315 ;
        RECT  355.015 0.17 355.785 0.94 ;
        RECT  355.015 0.17 355.275 12.9 ;
        RECT  355.525 0.17 355.785 12.9 ;
        RECT  354.515 190.585 354.715 191.315 ;
        RECT  355.015 190.585 355.215 191.315 ;
        RECT  355.51 190.585 355.71 191.315 ;
        RECT  356.035 0.52 356.295 5.815 ;
        RECT  356.89 0.52 357.15 5.16 ;
        RECT  356.89 4.9 357.67 5.16 ;
        RECT  357.41 4.9 357.67 6.64 ;
        RECT  356.33 190.585 356.53 191.315 ;
        RECT  356.825 190.585 357.025 191.315 ;
        RECT  357.325 190.585 357.525 191.315 ;
        RECT  357.825 190.585 358.025 191.315 ;
        RECT  358.32 190.585 358.52 191.315 ;
        RECT  359.14 190.585 359.34 191.315 ;
        RECT  359.635 190.585 359.835 191.315 ;
        RECT  360.135 190.585 360.335 191.315 ;
        RECT  360.29 0.52 360.55 2.335 ;
        RECT  360.635 190.585 360.835 191.315 ;
        RECT  360.8 0.52 361.06 14.11 ;
        RECT  361.13 190.585 361.33 191.315 ;
        RECT  362.175 0.17 362.945 0.94 ;
        RECT  362.685 0.17 362.945 8.7 ;
        RECT  362.175 0.17 362.435 12.9 ;
        RECT  361.665 0.52 361.925 2.485 ;
        RECT  361.95 190.585 362.15 191.315 ;
        RECT  363.195 0.17 363.965 0.43 ;
        RECT  363.705 0.17 363.965 10.48 ;
        RECT  363.195 0.17 363.455 10.99 ;
        RECT  362.445 190.585 362.645 191.315 ;
        RECT  362.945 190.585 363.145 191.315 ;
        RECT  363.445 190.585 363.645 191.315 ;
        RECT  363.94 190.585 364.14 191.315 ;
        RECT  365.235 0.17 366.005 0.43 ;
        RECT  365.235 0.17 365.495 11.5 ;
        RECT  365.745 0.17 366.005 11.5 ;
        RECT  364.76 190.585 364.96 191.315 ;
        RECT  365.255 190.585 365.455 191.315 ;
        RECT  366.255 0.17 367.025 0.94 ;
        RECT  366.255 0.17 366.515 12.9 ;
        RECT  366.765 0.17 367.025 12.9 ;
        RECT  365.755 190.585 365.955 191.315 ;
        RECT  366.255 190.585 366.455 191.315 ;
        RECT  366.75 190.585 366.95 191.315 ;
        RECT  367.275 0.52 367.535 5.815 ;
        RECT  368.13 0.52 368.39 5.16 ;
        RECT  368.13 4.9 368.91 5.16 ;
        RECT  368.65 4.9 368.91 6.64 ;
        RECT  367.57 190.585 367.77 191.315 ;
        RECT  368.065 190.585 368.265 191.315 ;
        RECT  368.565 190.585 368.765 191.315 ;
        RECT  369.065 190.585 369.265 191.315 ;
        RECT  369.56 190.585 369.76 191.315 ;
        RECT  370.38 190.585 370.58 191.315 ;
        RECT  370.875 190.585 371.075 191.315 ;
        RECT  371.375 190.585 371.575 191.315 ;
        RECT  371.53 0.52 371.79 2.335 ;
        RECT  371.875 190.585 372.075 191.315 ;
        RECT  372.04 0.52 372.3 14.11 ;
        RECT  372.37 190.585 372.57 191.315 ;
        RECT  373.415 0.17 374.185 0.94 ;
        RECT  373.925 0.17 374.185 8.7 ;
        RECT  373.415 0.17 373.675 12.9 ;
        RECT  372.905 0.52 373.165 2.485 ;
        RECT  373.19 190.585 373.39 191.315 ;
        RECT  374.435 0.17 375.205 0.43 ;
        RECT  374.945 0.17 375.205 10.48 ;
        RECT  374.435 0.17 374.695 10.99 ;
        RECT  373.685 190.585 373.885 191.315 ;
        RECT  374.185 190.585 374.385 191.315 ;
        RECT  374.685 190.585 374.885 191.315 ;
        RECT  375.18 190.585 375.38 191.315 ;
        RECT  376.475 0.17 377.245 0.43 ;
        RECT  376.475 0.17 376.735 11.5 ;
        RECT  376.985 0.17 377.245 11.5 ;
        RECT  376 190.585 376.2 191.315 ;
        RECT  376.495 190.585 376.695 191.315 ;
        RECT  377.495 0.17 378.265 0.94 ;
        RECT  377.495 0.17 377.755 12.9 ;
        RECT  378.005 0.17 378.265 12.9 ;
        RECT  376.995 190.585 377.195 191.315 ;
        RECT  377.495 190.585 377.695 191.315 ;
        RECT  377.99 190.585 378.19 191.315 ;
        RECT  378.515 0.52 378.775 5.815 ;
        RECT  379.37 0.52 379.63 5.16 ;
        RECT  379.37 4.9 380.15 5.16 ;
        RECT  379.89 4.9 380.15 6.64 ;
        RECT  378.81 190.585 379.01 191.315 ;
        RECT  379.305 190.585 379.505 191.315 ;
        RECT  379.805 190.585 380.005 191.315 ;
        RECT  380.305 190.585 380.505 191.315 ;
        RECT  380.8 190.585 381 191.315 ;
        RECT  381.62 190.585 381.82 191.315 ;
        RECT  382.115 190.585 382.315 191.315 ;
        RECT  382.615 190.585 382.815 191.315 ;
        RECT  382.77 0.52 383.03 2.335 ;
        RECT  383.115 190.585 383.315 191.315 ;
        RECT  383.28 0.52 383.54 14.11 ;
        RECT  383.61 190.585 383.81 191.315 ;
        RECT  384.655 0.17 385.425 0.94 ;
        RECT  385.165 0.17 385.425 8.7 ;
        RECT  384.655 0.17 384.915 12.9 ;
        RECT  384.145 0.52 384.405 2.485 ;
        RECT  384.43 190.585 384.63 191.315 ;
        RECT  385.675 0.17 386.445 0.43 ;
        RECT  386.185 0.17 386.445 10.48 ;
        RECT  385.675 0.17 385.935 10.99 ;
        RECT  384.925 190.585 385.125 191.315 ;
        RECT  385.425 190.585 385.625 191.315 ;
        RECT  385.925 190.585 386.125 191.315 ;
        RECT  386.42 190.585 386.62 191.315 ;
        RECT  387.715 0.17 388.485 0.43 ;
        RECT  387.715 0.17 387.975 11.5 ;
        RECT  388.225 0.17 388.485 11.5 ;
        RECT  387.24 190.585 387.44 191.315 ;
        RECT  387.735 190.585 387.935 191.315 ;
        RECT  388.735 0.17 389.505 0.94 ;
        RECT  388.735 0.17 388.995 12.9 ;
        RECT  389.245 0.17 389.505 12.9 ;
        RECT  388.235 190.585 388.435 191.315 ;
        RECT  388.735 190.585 388.935 191.315 ;
        RECT  389.23 190.585 389.43 191.315 ;
        RECT  389.755 0.52 390.015 5.815 ;
        RECT  390.61 0.52 390.87 5.16 ;
        RECT  390.61 4.9 391.39 5.16 ;
        RECT  391.13 4.9 391.39 6.64 ;
        RECT  390.05 190.585 390.25 191.315 ;
        RECT  390.545 190.585 390.745 191.315 ;
        RECT  391.045 190.585 391.245 191.315 ;
        RECT  391.545 190.585 391.745 191.315 ;
        RECT  392.04 190.585 392.24 191.315 ;
        RECT  392.86 190.585 393.06 191.315 ;
        RECT  393.355 190.585 393.555 191.315 ;
        RECT  393.855 190.585 394.055 191.315 ;
        RECT  394.01 0.52 394.27 2.335 ;
        RECT  394.355 190.585 394.555 191.315 ;
        RECT  394.52 0.52 394.78 14.11 ;
        RECT  394.85 190.585 395.05 191.315 ;
        RECT  395.895 0.17 396.665 0.94 ;
        RECT  396.405 0.17 396.665 8.7 ;
        RECT  395.895 0.17 396.155 12.9 ;
        RECT  395.385 0.52 395.645 2.485 ;
        RECT  395.67 190.585 395.87 191.315 ;
        RECT  396.915 0.17 397.685 0.43 ;
        RECT  397.425 0.17 397.685 10.48 ;
        RECT  396.915 0.17 397.175 10.99 ;
        RECT  396.165 190.585 396.365 191.315 ;
        RECT  396.665 190.585 396.865 191.315 ;
        RECT  397.165 190.585 397.365 191.315 ;
        RECT  397.66 190.585 397.86 191.315 ;
        RECT  398.955 0.17 399.725 0.43 ;
        RECT  398.955 0.17 399.215 11.5 ;
        RECT  399.465 0.17 399.725 11.5 ;
        RECT  398.48 190.585 398.68 191.315 ;
        RECT  398.975 190.585 399.175 191.315 ;
        RECT  399.975 0.17 400.745 0.94 ;
        RECT  399.975 0.17 400.235 12.9 ;
        RECT  400.485 0.17 400.745 12.9 ;
        RECT  399.475 190.585 399.675 191.315 ;
        RECT  399.975 190.585 400.175 191.315 ;
        RECT  400.47 190.585 400.67 191.315 ;
        RECT  400.995 0.52 401.255 5.815 ;
        RECT  401.85 0.52 402.11 5.16 ;
        RECT  401.85 4.9 402.63 5.16 ;
        RECT  402.37 4.9 402.63 6.64 ;
        RECT  401.29 190.585 401.49 191.315 ;
        RECT  401.785 190.585 401.985 191.315 ;
        RECT  402.285 190.585 402.485 191.315 ;
        RECT  402.785 190.585 402.985 191.315 ;
        RECT  403.28 190.585 403.48 191.315 ;
        RECT  404.1 190.585 404.3 191.315 ;
        RECT  404.595 190.585 404.795 191.315 ;
        RECT  405.095 190.585 405.295 191.315 ;
        RECT  405.25 0.52 405.51 2.335 ;
        RECT  405.595 190.585 405.795 191.315 ;
        RECT  405.76 0.52 406.02 14.11 ;
        RECT  406.09 190.585 406.29 191.315 ;
        RECT  407.135 0.17 407.905 0.94 ;
        RECT  407.645 0.17 407.905 8.7 ;
        RECT  407.135 0.17 407.395 12.9 ;
        RECT  406.625 0.52 406.885 2.485 ;
        RECT  406.91 190.585 407.11 191.315 ;
        RECT  408.155 0.17 408.925 0.43 ;
        RECT  408.665 0.17 408.925 10.48 ;
        RECT  408.155 0.17 408.415 10.99 ;
        RECT  407.405 190.585 407.605 191.315 ;
        RECT  407.905 190.585 408.105 191.315 ;
        RECT  408.405 190.585 408.605 191.315 ;
        RECT  408.9 190.585 409.1 191.315 ;
        RECT  410.195 0.17 410.965 0.43 ;
        RECT  410.195 0.17 410.455 11.5 ;
        RECT  410.705 0.17 410.965 11.5 ;
        RECT  409.72 190.585 409.92 191.315 ;
        RECT  410.215 190.585 410.415 191.315 ;
        RECT  411.215 0.17 411.985 0.94 ;
        RECT  411.215 0.17 411.475 12.9 ;
        RECT  411.725 0.17 411.985 12.9 ;
        RECT  410.715 190.585 410.915 191.315 ;
        RECT  411.215 190.585 411.415 191.315 ;
        RECT  411.71 190.585 411.91 191.315 ;
        RECT  412.235 0.52 412.495 5.815 ;
        RECT  413.09 0.52 413.35 5.16 ;
        RECT  413.09 4.9 413.87 5.16 ;
        RECT  413.61 4.9 413.87 6.64 ;
        RECT  412.53 190.585 412.73 191.315 ;
        RECT  413.025 190.585 413.225 191.315 ;
        RECT  413.525 190.585 413.725 191.315 ;
        RECT  414.025 190.585 414.225 191.315 ;
        RECT  414.52 190.585 414.72 191.315 ;
        RECT  415.34 190.585 415.54 191.315 ;
        RECT  416.335 45.465 416.535 191.315 ;
        RECT  249.785 0 254.615 191.34 ;
        RECT  261.025 0 265.855 191.34 ;
        RECT  272.265 0 277.095 191.34 ;
        RECT  283.505 0 288.335 191.34 ;
        RECT  294.745 0 299.575 191.34 ;
        RECT  305.985 0 310.815 191.34 ;
        RECT  317.225 0 322.055 191.34 ;
        RECT  328.465 0 333.295 191.34 ;
        RECT  339.705 0 344.535 191.34 ;
        RECT  350.945 0 355.775 191.34 ;
        RECT  362.185 0 367.015 191.34 ;
        RECT  373.425 0 378.255 191.34 ;
        RECT  384.665 0 389.495 191.34 ;
        RECT  395.905 0 400.735 191.34 ;
        RECT  407.145 0 411.975 191.34 ;
        RECT  201.98 0 202.22 191.34 ;
        RECT  203.51 0 203.75 191.34 ;
        RECT  206.57 0 206.81 191.34 ;
        RECT  208.1 0 208.34 191.34 ;
        RECT  215.23 0 222.11 191.34 ;
        RECT  223.4 0 224.15 191.34 ;
        RECT  0 0 3.03 191.34 ;
        RECT  4.655 0.17 9.505 191.34 ;
        RECT  11.65 0 14.27 191.34 ;
        RECT  15.895 0.17 20.745 191.34 ;
        RECT  22.89 0 25.51 191.34 ;
        RECT  27.135 0.17 31.985 191.34 ;
        RECT  34.13 0 36.75 191.34 ;
        RECT  38.375 0.17 43.225 191.34 ;
        RECT  45.37 0 47.99 191.34 ;
        RECT  49.615 0.17 54.465 191.34 ;
        RECT  56.61 0 59.23 191.34 ;
        RECT  60.855 0.17 65.705 191.34 ;
        RECT  67.85 0 70.47 191.34 ;
        RECT  72.095 0.17 76.945 191.34 ;
        RECT  79.09 0 81.71 191.34 ;
        RECT  83.335 0.17 88.185 191.34 ;
        RECT  90.33 0 92.95 191.34 ;
        RECT  94.575 0.17 99.425 191.34 ;
        RECT  101.57 0 104.19 191.34 ;
        RECT  105.815 0.17 110.665 191.34 ;
        RECT  112.81 0 115.43 191.34 ;
        RECT  117.055 0.17 121.905 191.34 ;
        RECT  124.05 0 126.67 191.34 ;
        RECT  128.295 0.17 133.145 191.34 ;
        RECT  135.29 0 137.91 191.34 ;
        RECT  139.535 0.17 144.385 191.34 ;
        RECT  146.53 0 149.15 191.34 ;
        RECT  150.775 0.17 155.625 191.34 ;
        RECT  157.77 0 160.39 191.34 ;
        RECT  162.015 0.17 166.865 191.34 ;
        RECT  169.01 0 171.63 191.34 ;
        RECT  173.255 0.17 178.105 191.34 ;
        RECT  180.25 0 192.03 191.34 ;
        RECT  194.32 0.17 200.7 191.34 ;
        RECT  201.97 0.3 202.23 191.34 ;
        RECT  203.5 0.3 203.76 191.34 ;
        RECT  206.56 0.3 206.82 191.34 ;
        RECT  208.09 0.3 208.35 191.34 ;
        RECT  209.63 0.17 210.9 191.34 ;
        RECT  209.62 0.3 210.9 191.34 ;
        RECT  215.23 0.3 222.12 191.34 ;
        RECT  223.39 0.3 224.16 191.34 ;
        RECT  224.93 0 236.39 191.34 ;
        RECT  224.92 0.17 236.39 191.34 ;
        RECT  238.535 0.17 243.385 191.34 ;
        RECT  245.01 0 247.63 191.34 ;
        RECT  249.775 0.17 254.625 191.34 ;
        RECT  256.25 0 258.87 191.34 ;
        RECT  261.015 0.17 265.865 191.34 ;
        RECT  267.49 0 270.11 191.34 ;
        RECT  272.255 0.17 277.105 191.34 ;
        RECT  278.73 0 281.35 191.34 ;
        RECT  283.495 0.17 288.345 191.34 ;
        RECT  289.97 0 292.59 191.34 ;
        RECT  294.735 0.17 299.585 191.34 ;
        RECT  301.21 0 303.83 191.34 ;
        RECT  305.975 0.17 310.825 191.34 ;
        RECT  312.45 0 315.07 191.34 ;
        RECT  317.215 0.17 322.065 191.34 ;
        RECT  323.69 0 326.31 191.34 ;
        RECT  328.455 0.17 333.305 191.34 ;
        RECT  334.93 0 337.55 191.34 ;
        RECT  339.695 0.17 344.545 191.34 ;
        RECT  346.17 0 348.79 191.34 ;
        RECT  350.935 0.17 355.785 191.34 ;
        RECT  357.41 0 360.03 191.34 ;
        RECT  362.175 0.17 367.025 191.34 ;
        RECT  368.65 0 371.27 191.34 ;
        RECT  373.415 0.17 378.265 191.34 ;
        RECT  379.89 0 382.51 191.34 ;
        RECT  384.655 0.17 389.505 191.34 ;
        RECT  391.13 0 393.75 191.34 ;
        RECT  395.895 0.17 400.745 191.34 ;
        RECT  402.37 0 404.99 191.34 ;
        RECT  407.135 0.17 411.985 191.34 ;
        RECT  413.61 0 416.64 191.34 ;
        RECT  0 0.52 416.64 191.34 ;
        RECT  4.665 0 9.495 191.34 ;
        RECT  15.905 0 20.735 191.34 ;
        RECT  27.145 0 31.975 191.34 ;
        RECT  38.385 0 43.215 191.34 ;
        RECT  49.625 0 54.455 191.34 ;
        RECT  60.865 0 65.695 191.34 ;
        RECT  72.105 0 76.935 191.34 ;
        RECT  83.345 0 88.175 191.34 ;
        RECT  94.585 0 99.415 191.34 ;
        RECT  105.825 0 110.655 191.34 ;
        RECT  117.065 0 121.895 191.34 ;
        RECT  128.305 0 133.135 191.34 ;
        RECT  139.545 0 144.375 191.34 ;
        RECT  150.785 0 155.615 191.34 ;
        RECT  162.025 0 166.855 191.34 ;
        RECT  173.265 0 178.095 191.34 ;
        RECT  194.32 0 200.69 191.34 ;
        RECT  209.63 0 210.89 191.34 ;
        RECT  238.545 0 243.375 191.34 ;
      LAYER Metal3 ;
        RECT  0 0 416.64 191.34 ;
      LAYER Metal4 ;
        RECT  0 39.085 9.62 45.205 ;
        RECT  0 0 4 191.34 ;
        RECT  7.33 0 9.62 191.34 ;
        RECT  12.95 39.085 20.86 45.205 ;
        RECT  12.95 0 15.24 191.34 ;
        RECT  18.57 0 20.86 191.34 ;
        RECT  24.19 39.085 32.1 45.205 ;
        RECT  24.19 0 26.48 191.34 ;
        RECT  29.81 0 32.1 191.34 ;
        RECT  35.43 39.085 43.34 45.205 ;
        RECT  35.43 0 37.72 191.34 ;
        RECT  41.05 0 43.34 191.34 ;
        RECT  46.67 39.085 54.58 45.205 ;
        RECT  46.67 0 48.96 191.34 ;
        RECT  52.29 0 54.58 191.34 ;
        RECT  57.91 39.085 65.82 45.205 ;
        RECT  57.91 0 60.2 191.34 ;
        RECT  63.53 0 65.82 191.34 ;
        RECT  69.15 39.085 77.06 45.205 ;
        RECT  69.15 0 71.44 191.34 ;
        RECT  74.77 0 77.06 191.34 ;
        RECT  80.39 39.085 88.3 45.205 ;
        RECT  80.39 0 82.68 191.34 ;
        RECT  86.01 0 88.3 191.34 ;
        RECT  91.63 39.085 99.54 45.205 ;
        RECT  91.63 0 93.92 191.34 ;
        RECT  97.25 0 99.54 191.34 ;
        RECT  102.87 39.085 110.78 45.205 ;
        RECT  102.87 0 105.16 191.34 ;
        RECT  108.49 0 110.78 191.34 ;
        RECT  114.11 39.085 122.02 45.205 ;
        RECT  114.11 0 116.4 191.34 ;
        RECT  119.73 0 122.02 191.34 ;
        RECT  125.35 39.085 133.26 45.205 ;
        RECT  125.35 0 127.64 191.34 ;
        RECT  130.97 0 133.26 191.34 ;
        RECT  136.59 39.085 144.5 45.205 ;
        RECT  136.59 0 138.88 191.34 ;
        RECT  142.21 0 144.5 191.34 ;
        RECT  147.83 39.085 155.74 45.205 ;
        RECT  147.83 0 150.12 191.34 ;
        RECT  153.45 0 155.74 191.34 ;
        RECT  159.07 39.085 166.98 45.205 ;
        RECT  159.07 0 161.36 191.34 ;
        RECT  164.69 0 166.98 191.34 ;
        RECT  170.31 39.085 178.22 45.205 ;
        RECT  170.31 0 172.6 191.34 ;
        RECT  175.93 0 178.22 191.34 ;
        RECT  181.55 0 188.63 191.34 ;
        RECT  191.96 0 193.78 191.34 ;
        RECT  197.11 0 198.93 191.34 ;
        RECT  202.26 0 204.08 191.34 ;
        RECT  207.41 0 209.23 191.34 ;
        RECT  212.56 0 214.38 191.34 ;
        RECT  238.42 39.085 246.33 45.205 ;
        RECT  238.42 0 240.71 191.34 ;
        RECT  244.04 0 246.33 191.34 ;
        RECT  249.66 39.085 257.57 45.205 ;
        RECT  249.66 0 251.95 191.34 ;
        RECT  255.28 0 257.57 191.34 ;
        RECT  260.9 39.085 268.81 45.205 ;
        RECT  260.9 0 263.19 191.34 ;
        RECT  266.52 0 268.81 191.34 ;
        RECT  272.14 39.085 280.05 45.205 ;
        RECT  272.14 0 274.43 191.34 ;
        RECT  277.76 0 280.05 191.34 ;
        RECT  283.38 39.085 291.29 45.205 ;
        RECT  283.38 0 285.67 191.34 ;
        RECT  289 0 291.29 191.34 ;
        RECT  294.62 39.085 302.53 45.205 ;
        RECT  294.62 0 296.91 191.34 ;
        RECT  300.24 0 302.53 191.34 ;
        RECT  305.86 39.085 313.77 45.205 ;
        RECT  305.86 0 308.15 191.34 ;
        RECT  311.48 0 313.77 191.34 ;
        RECT  317.1 39.085 325.01 45.205 ;
        RECT  317.1 0 319.39 191.34 ;
        RECT  322.72 0 325.01 191.34 ;
        RECT  328.34 39.085 336.25 45.205 ;
        RECT  328.34 0 330.63 191.34 ;
        RECT  333.96 0 336.25 191.34 ;
        RECT  339.58 39.085 347.49 45.205 ;
        RECT  339.58 0 341.87 191.34 ;
        RECT  345.2 0 347.49 191.34 ;
        RECT  350.82 39.085 358.73 45.205 ;
        RECT  350.82 0 353.11 191.34 ;
        RECT  356.44 0 358.73 191.34 ;
        RECT  362.06 39.085 369.97 45.205 ;
        RECT  362.06 0 364.35 191.34 ;
        RECT  367.68 0 369.97 191.34 ;
        RECT  373.3 39.085 381.21 45.205 ;
        RECT  373.3 0 375.59 191.34 ;
        RECT  378.92 0 381.21 191.34 ;
        RECT  384.54 39.085 392.45 45.205 ;
        RECT  384.54 0 386.83 191.34 ;
        RECT  390.16 0 392.45 191.34 ;
        RECT  395.78 39.085 403.69 45.205 ;
        RECT  395.78 0 398.07 191.34 ;
        RECT  401.4 0 403.69 191.34 ;
        RECT  407.02 39.085 416.64 45.205 ;
        RECT  407.02 0 409.31 191.34 ;
        RECT  412.64 0 416.64 191.34 ;
        RECT  217.71 0 219.53 191.34 ;
        RECT  222.86 0 224.68 191.34 ;
        RECT  228.01 0 235.09 191.34 ;
    END
END RM_IHPSG13_1P_512x32_c2_bm_bist
END LIBRARY
