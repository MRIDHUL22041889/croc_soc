VERSION 5.7 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "|" ;

PROPERTYDEFINITIONS
END PROPERTYDEFINITIONS


MACRO bondpad_70x70
    CLASS COVER ;
    SIZE 70 BY 70 ;
    SYMMETRY X Y R90 ;
    SITE sg13g2_ioSite ;
    PIN pad
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal2 ;
              RECT  0 0 70 70 ;
            LAYER Metal3 ;
              RECT  0 0 70 70 ;
            LAYER Metal4 ;
              RECT  0 0 70 70 ;
            LAYER Metal5 ;
              RECT  0 0 70 70 ;
            LAYER TopMetal1 ;
              RECT  0 0 70 70 ;
            LAYER TopMetal2 ;
              RECT  0 0 70 70 ;
        END
    END pad
    OBS
      LAYER Metal1 ;
        RECT  0 0 70 70 ;
      LAYER Metal2 ;
        RECT  0 0 70 70 ;
      LAYER Metal3 ;
        RECT  0 0 70 70 ;
      LAYER Metal4 ;
        RECT  0 0 70 70 ;
      LAYER Metal5 ;
        RECT  0 0 70 70 ;
      LAYER TopMetal1 ;
        RECT  0 0 70 70 ;
      LAYER TopMetal2 ;
        RECT  0 0 70 70 ;
    END
END bondpad_70x70
END LIBRARY
