VERSION 5.7 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

PROPERTYDEFINITIONS
END PROPERTYDEFINITIONS


MACRO RM_IHPSG13_1P_512x64_c2_bm_bist
    CLASS BLOCK ;
    SIZE 784.48 BY 191.34 ;
    SYMMETRY X Y R90 ;
    PIN A_DIN[32]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  432.49 0 432.75 0.26 ;
        END
    END A_DIN[32]
    PIN A_DIN[31]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  351.73 0 351.99 0.26 ;
        END
    END A_DIN[31]
    PIN A_BIST_DIN[32]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  431.635 0 431.895 0.26 ;
        END
    END A_BIST_DIN[32]
    PIN A_BIST_DIN[31]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  352.585 0 352.845 0.26 ;
        END
    END A_BIST_DIN[31]
    PIN A_BM[32]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  424.65 0 424.91 0.26 ;
        END
    END A_BM[32]
    PIN A_BM[31]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  359.57 0 359.83 0.26 ;
        END
    END A_BM[31]
    PIN A_BIST_BM[32]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  426.025 0 426.285 0.26 ;
        END
    END A_BIST_BM[32]
    PIN A_BIST_BM[31]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  358.195 0 358.455 0.26 ;
        END
    END A_BIST_BM[31]
    PIN A_DOUT[32]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  425.16 0 425.42 0.26 ;
        END
    END A_DOUT[32]
    PIN A_DOUT[31]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  359.06 0 359.32 0.26 ;
        END
    END A_DOUT[31]
    PIN VSS!
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal4 ;
              RECT  771.79 0 774.6 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  760.55 0 763.36 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  749.31 0 752.12 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  738.07 0 740.88 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  726.83 0 729.64 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  715.59 0 718.4 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  704.35 0 707.16 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  693.11 0 695.92 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  681.87 0 684.68 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  670.63 0 673.44 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  659.39 0 662.2 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  648.15 0 650.96 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  636.91 0 639.72 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  625.67 0 628.48 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  614.43 0 617.24 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  603.19 0 606 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  591.95 0 594.76 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  580.71 0 583.52 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  569.47 0 572.28 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  558.23 0 561.04 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  546.99 0 549.8 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  535.75 0 538.56 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  524.51 0 527.32 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  513.27 0 516.08 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  502.03 0 504.84 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  490.79 0 493.6 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  479.55 0 482.36 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  468.31 0 471.12 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  457.07 0 459.88 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  445.83 0 448.64 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  434.59 0 437.4 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  423.35 0 426.16 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  408.86 0 411.67 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  398.56 0 401.37 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  383.11 0 385.92 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  372.81 0 375.62 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  358.32 0 361.13 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  347.08 0 349.89 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  335.84 0 338.65 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  324.6 0 327.41 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  313.36 0 316.17 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  302.12 0 304.93 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  290.88 0 293.69 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  279.64 0 282.45 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  268.4 0 271.21 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  257.16 0 259.97 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  245.92 0 248.73 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  234.68 0 237.49 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  223.44 0 226.25 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  212.2 0 215.01 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  200.96 0 203.77 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  189.72 0 192.53 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  178.48 0 181.29 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  167.24 0 170.05 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  156 0 158.81 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  144.76 0 147.57 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  133.52 0 136.33 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  122.28 0 125.09 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  111.04 0 113.85 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  99.8 0 102.61 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  88.56 0 91.37 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  77.32 0 80.13 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  66.08 0 68.89 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  54.84 0 57.65 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  43.6 0 46.41 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  32.36 0 35.17 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  21.12 0 23.93 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  9.88 0 12.69 191.34 ;
        END
    END VSS!
    PIN VDD!
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal4 ;
              RECT  777.41 0 780.22 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  766.17 0 768.98 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  754.93 0 757.74 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  743.69 0 746.5 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  732.45 0 735.26 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  721.21 0 724.02 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  709.97 0 712.78 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  698.73 0 701.54 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  687.49 0 690.3 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  676.25 0 679.06 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  665.01 0 667.82 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  653.77 0 656.58 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  642.53 0 645.34 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  631.29 0 634.1 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  620.05 0 622.86 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  608.81 0 611.62 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  597.57 0 600.38 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  586.33 0 589.14 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  575.09 0 577.9 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  563.85 0 566.66 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  552.61 0 555.42 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  541.37 0 544.18 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  530.13 0 532.94 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  518.89 0 521.7 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  507.65 0 510.46 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  496.41 0 499.22 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  485.17 0 487.98 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  473.93 0 476.74 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  462.69 0 465.5 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  451.45 0 454.26 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  440.21 0 443.02 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  428.97 0 431.78 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  403.71 0 406.52 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  393.41 0 396.22 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  388.26 0 391.07 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  377.96 0 380.77 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  352.7 0 355.51 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  341.46 0 344.27 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  330.22 0 333.03 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  318.98 0 321.79 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  307.74 0 310.55 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  296.5 0 299.31 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  285.26 0 288.07 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  274.02 0 276.83 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  262.78 0 265.59 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  251.54 0 254.35 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  240.3 0 243.11 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  229.06 0 231.87 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  217.82 0 220.63 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  206.58 0 209.39 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  195.34 0 198.15 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  184.1 0 186.91 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  172.86 0 175.67 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  161.62 0 164.43 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  150.38 0 153.19 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  139.14 0 141.95 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  127.9 0 130.71 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  116.66 0 119.47 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  105.42 0 108.23 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  94.18 0 96.99 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  82.94 0 85.75 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  71.7 0 74.51 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  60.46 0 63.27 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  49.22 0 52.03 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  37.98 0 40.79 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  26.74 0 29.55 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  15.5 0 18.31 38.825 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  4.26 0 7.07 38.825 ;
        END
    END VDD!
    PIN VDDARRAY!
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal4 ;
              RECT  777.41 45.465 780.22 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  766.17 45.465 768.98 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  754.93 45.465 757.74 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  743.69 45.465 746.5 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  732.45 45.465 735.26 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  721.21 45.465 724.02 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  709.97 45.465 712.78 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  698.73 45.465 701.54 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  687.49 45.465 690.3 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  676.25 45.465 679.06 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  665.01 45.465 667.82 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  653.77 45.465 656.58 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  642.53 45.465 645.34 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  631.29 45.465 634.1 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  620.05 45.465 622.86 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  608.81 45.465 611.62 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  597.57 45.465 600.38 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  586.33 45.465 589.14 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  575.09 45.465 577.9 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  563.85 45.465 566.66 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  552.61 45.465 555.42 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  541.37 45.465 544.18 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  530.13 45.465 532.94 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  518.89 45.465 521.7 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  507.65 45.465 510.46 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  496.41 45.465 499.22 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  485.17 45.465 487.98 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  473.93 45.465 476.74 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  462.69 45.465 465.5 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  451.45 45.465 454.26 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  440.21 45.465 443.02 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  428.97 45.465 431.78 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  352.7 45.465 355.51 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  341.46 45.465 344.27 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  330.22 45.465 333.03 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  318.98 45.465 321.79 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  307.74 45.465 310.55 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  296.5 45.465 299.31 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  285.26 45.465 288.07 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  274.02 45.465 276.83 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  262.78 45.465 265.59 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  251.54 45.465 254.35 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  240.3 45.465 243.11 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  229.06 45.465 231.87 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  217.82 45.465 220.63 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  206.58 45.465 209.39 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  195.34 45.465 198.15 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  184.1 45.465 186.91 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  172.86 45.465 175.67 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  161.62 45.465 164.43 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  150.38 45.465 153.19 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  139.14 45.465 141.95 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  127.9 45.465 130.71 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  116.66 45.465 119.47 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  105.42 45.465 108.23 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  94.18 45.465 96.99 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  82.94 45.465 85.75 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  71.7 45.465 74.51 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  60.46 45.465 63.27 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  49.22 45.465 52.03 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  37.98 45.465 40.79 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  26.74 45.465 29.55 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  15.5 45.465 18.31 191.34 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  4.26 45.465 7.07 191.34 ;
        END
    END VDDARRAY!
    PIN A_DIN[33]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  443.73 0 443.99 0.26 ;
        END
    END A_DIN[33]
    PIN A_DIN[30]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  340.49 0 340.75 0.26 ;
        END
    END A_DIN[30]
    PIN A_BIST_DIN[33]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  442.875 0 443.135 0.26 ;
        END
    END A_BIST_DIN[33]
    PIN A_BIST_DIN[30]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  341.345 0 341.605 0.26 ;
        END
    END A_BIST_DIN[30]
    PIN A_BM[33]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  435.89 0 436.15 0.26 ;
        END
    END A_BM[33]
    PIN A_BM[30]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  348.33 0 348.59 0.26 ;
        END
    END A_BM[30]
    PIN A_BIST_BM[33]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  437.265 0 437.525 0.26 ;
        END
    END A_BIST_BM[33]
    PIN A_BIST_BM[30]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  346.955 0 347.215 0.26 ;
        END
    END A_BIST_BM[30]
    PIN A_DOUT[33]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  436.4 0 436.66 0.26 ;
        END
    END A_DOUT[33]
    PIN A_DOUT[30]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  347.82 0 348.08 0.26 ;
        END
    END A_DOUT[30]
    PIN A_DIN[34]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  454.97 0 455.23 0.26 ;
        END
    END A_DIN[34]
    PIN A_DIN[29]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  329.25 0 329.51 0.26 ;
        END
    END A_DIN[29]
    PIN A_BIST_DIN[34]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  454.115 0 454.375 0.26 ;
        END
    END A_BIST_DIN[34]
    PIN A_BIST_DIN[29]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  330.105 0 330.365 0.26 ;
        END
    END A_BIST_DIN[29]
    PIN A_BM[34]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  447.13 0 447.39 0.26 ;
        END
    END A_BM[34]
    PIN A_BM[29]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  337.09 0 337.35 0.26 ;
        END
    END A_BM[29]
    PIN A_BIST_BM[34]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  448.505 0 448.765 0.26 ;
        END
    END A_BIST_BM[34]
    PIN A_BIST_BM[29]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  335.715 0 335.975 0.26 ;
        END
    END A_BIST_BM[29]
    PIN A_DOUT[34]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  447.64 0 447.9 0.26 ;
        END
    END A_DOUT[34]
    PIN A_DOUT[29]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  336.58 0 336.84 0.26 ;
        END
    END A_DOUT[29]
    PIN A_DIN[35]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  466.21 0 466.47 0.26 ;
        END
    END A_DIN[35]
    PIN A_DIN[28]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  318.01 0 318.27 0.26 ;
        END
    END A_DIN[28]
    PIN A_BIST_DIN[35]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  465.355 0 465.615 0.26 ;
        END
    END A_BIST_DIN[35]
    PIN A_BIST_DIN[28]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  318.865 0 319.125 0.26 ;
        END
    END A_BIST_DIN[28]
    PIN A_BM[35]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  458.37 0 458.63 0.26 ;
        END
    END A_BM[35]
    PIN A_BM[28]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  325.85 0 326.11 0.26 ;
        END
    END A_BM[28]
    PIN A_BIST_BM[35]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  459.745 0 460.005 0.26 ;
        END
    END A_BIST_BM[35]
    PIN A_BIST_BM[28]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  324.475 0 324.735 0.26 ;
        END
    END A_BIST_BM[28]
    PIN A_DOUT[35]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  458.88 0 459.14 0.26 ;
        END
    END A_DOUT[35]
    PIN A_DOUT[28]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  325.34 0 325.6 0.26 ;
        END
    END A_DOUT[28]
    PIN A_DIN[36]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  477.45 0 477.71 0.26 ;
        END
    END A_DIN[36]
    PIN A_DIN[27]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  306.77 0 307.03 0.26 ;
        END
    END A_DIN[27]
    PIN A_BIST_DIN[36]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  476.595 0 476.855 0.26 ;
        END
    END A_BIST_DIN[36]
    PIN A_BIST_DIN[27]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  307.625 0 307.885 0.26 ;
        END
    END A_BIST_DIN[27]
    PIN A_BM[36]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  469.61 0 469.87 0.26 ;
        END
    END A_BM[36]
    PIN A_BM[27]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  314.61 0 314.87 0.26 ;
        END
    END A_BM[27]
    PIN A_BIST_BM[36]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  470.985 0 471.245 0.26 ;
        END
    END A_BIST_BM[36]
    PIN A_BIST_BM[27]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  313.235 0 313.495 0.26 ;
        END
    END A_BIST_BM[27]
    PIN A_DOUT[36]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  470.12 0 470.38 0.26 ;
        END
    END A_DOUT[36]
    PIN A_DOUT[27]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  314.1 0 314.36 0.26 ;
        END
    END A_DOUT[27]
    PIN A_DIN[37]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  488.69 0 488.95 0.26 ;
        END
    END A_DIN[37]
    PIN A_DIN[26]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  295.53 0 295.79 0.26 ;
        END
    END A_DIN[26]
    PIN A_BIST_DIN[37]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  487.835 0 488.095 0.26 ;
        END
    END A_BIST_DIN[37]
    PIN A_BIST_DIN[26]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  296.385 0 296.645 0.26 ;
        END
    END A_BIST_DIN[26]
    PIN A_BM[37]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  480.85 0 481.11 0.26 ;
        END
    END A_BM[37]
    PIN A_BM[26]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  303.37 0 303.63 0.26 ;
        END
    END A_BM[26]
    PIN A_BIST_BM[37]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  482.225 0 482.485 0.26 ;
        END
    END A_BIST_BM[37]
    PIN A_BIST_BM[26]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  301.995 0 302.255 0.26 ;
        END
    END A_BIST_BM[26]
    PIN A_DOUT[37]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  481.36 0 481.62 0.26 ;
        END
    END A_DOUT[37]
    PIN A_DOUT[26]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  302.86 0 303.12 0.26 ;
        END
    END A_DOUT[26]
    PIN A_DIN[38]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  499.93 0 500.19 0.26 ;
        END
    END A_DIN[38]
    PIN A_DIN[25]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  284.29 0 284.55 0.26 ;
        END
    END A_DIN[25]
    PIN A_BIST_DIN[38]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  499.075 0 499.335 0.26 ;
        END
    END A_BIST_DIN[38]
    PIN A_BIST_DIN[25]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  285.145 0 285.405 0.26 ;
        END
    END A_BIST_DIN[25]
    PIN A_BM[38]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  492.09 0 492.35 0.26 ;
        END
    END A_BM[38]
    PIN A_BM[25]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  292.13 0 292.39 0.26 ;
        END
    END A_BM[25]
    PIN A_BIST_BM[38]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  493.465 0 493.725 0.26 ;
        END
    END A_BIST_BM[38]
    PIN A_BIST_BM[25]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  290.755 0 291.015 0.26 ;
        END
    END A_BIST_BM[25]
    PIN A_DOUT[38]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  492.6 0 492.86 0.26 ;
        END
    END A_DOUT[38]
    PIN A_DOUT[25]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  291.62 0 291.88 0.26 ;
        END
    END A_DOUT[25]
    PIN A_DIN[39]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  511.17 0 511.43 0.26 ;
        END
    END A_DIN[39]
    PIN A_DIN[24]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  273.05 0 273.31 0.26 ;
        END
    END A_DIN[24]
    PIN A_BIST_DIN[39]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  510.315 0 510.575 0.26 ;
        END
    END A_BIST_DIN[39]
    PIN A_BIST_DIN[24]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  273.905 0 274.165 0.26 ;
        END
    END A_BIST_DIN[24]
    PIN A_BM[39]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  503.33 0 503.59 0.26 ;
        END
    END A_BM[39]
    PIN A_BM[24]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  280.89 0 281.15 0.26 ;
        END
    END A_BM[24]
    PIN A_BIST_BM[39]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  504.705 0 504.965 0.26 ;
        END
    END A_BIST_BM[39]
    PIN A_BIST_BM[24]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  279.515 0 279.775 0.26 ;
        END
    END A_BIST_BM[24]
    PIN A_DOUT[39]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  503.84 0 504.1 0.26 ;
        END
    END A_DOUT[39]
    PIN A_DOUT[24]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  280.38 0 280.64 0.26 ;
        END
    END A_DOUT[24]
    PIN A_DIN[40]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  522.41 0 522.67 0.26 ;
        END
    END A_DIN[40]
    PIN A_DIN[23]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  261.81 0 262.07 0.26 ;
        END
    END A_DIN[23]
    PIN A_BIST_DIN[40]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  521.555 0 521.815 0.26 ;
        END
    END A_BIST_DIN[40]
    PIN A_BIST_DIN[23]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  262.665 0 262.925 0.26 ;
        END
    END A_BIST_DIN[23]
    PIN A_BM[40]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  514.57 0 514.83 0.26 ;
        END
    END A_BM[40]
    PIN A_BM[23]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  269.65 0 269.91 0.26 ;
        END
    END A_BM[23]
    PIN A_BIST_BM[40]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  515.945 0 516.205 0.26 ;
        END
    END A_BIST_BM[40]
    PIN A_BIST_BM[23]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  268.275 0 268.535 0.26 ;
        END
    END A_BIST_BM[23]
    PIN A_DOUT[40]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  515.08 0 515.34 0.26 ;
        END
    END A_DOUT[40]
    PIN A_DOUT[23]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  269.14 0 269.4 0.26 ;
        END
    END A_DOUT[23]
    PIN A_DIN[41]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  533.65 0 533.91 0.26 ;
        END
    END A_DIN[41]
    PIN A_DIN[22]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  250.57 0 250.83 0.26 ;
        END
    END A_DIN[22]
    PIN A_BIST_DIN[41]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  532.795 0 533.055 0.26 ;
        END
    END A_BIST_DIN[41]
    PIN A_BIST_DIN[22]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  251.425 0 251.685 0.26 ;
        END
    END A_BIST_DIN[22]
    PIN A_BM[41]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  525.81 0 526.07 0.26 ;
        END
    END A_BM[41]
    PIN A_BM[22]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  258.41 0 258.67 0.26 ;
        END
    END A_BM[22]
    PIN A_BIST_BM[41]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  527.185 0 527.445 0.26 ;
        END
    END A_BIST_BM[41]
    PIN A_BIST_BM[22]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  257.035 0 257.295 0.26 ;
        END
    END A_BIST_BM[22]
    PIN A_DOUT[41]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  526.32 0 526.58 0.26 ;
        END
    END A_DOUT[41]
    PIN A_DOUT[22]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  257.9 0 258.16 0.26 ;
        END
    END A_DOUT[22]
    PIN A_DIN[42]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  544.89 0 545.15 0.26 ;
        END
    END A_DIN[42]
    PIN A_DIN[21]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  239.33 0 239.59 0.26 ;
        END
    END A_DIN[21]
    PIN A_BIST_DIN[42]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  544.035 0 544.295 0.26 ;
        END
    END A_BIST_DIN[42]
    PIN A_BIST_DIN[21]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  240.185 0 240.445 0.26 ;
        END
    END A_BIST_DIN[21]
    PIN A_BM[42]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  537.05 0 537.31 0.26 ;
        END
    END A_BM[42]
    PIN A_BM[21]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  247.17 0 247.43 0.26 ;
        END
    END A_BM[21]
    PIN A_BIST_BM[42]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  538.425 0 538.685 0.26 ;
        END
    END A_BIST_BM[42]
    PIN A_BIST_BM[21]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  245.795 0 246.055 0.26 ;
        END
    END A_BIST_BM[21]
    PIN A_DOUT[42]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  537.56 0 537.82 0.26 ;
        END
    END A_DOUT[42]
    PIN A_DOUT[21]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  246.66 0 246.92 0.26 ;
        END
    END A_DOUT[21]
    PIN A_DIN[43]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  556.13 0 556.39 0.26 ;
        END
    END A_DIN[43]
    PIN A_DIN[20]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  228.09 0 228.35 0.26 ;
        END
    END A_DIN[20]
    PIN A_BIST_DIN[43]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  555.275 0 555.535 0.26 ;
        END
    END A_BIST_DIN[43]
    PIN A_BIST_DIN[20]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  228.945 0 229.205 0.26 ;
        END
    END A_BIST_DIN[20]
    PIN A_BM[43]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  548.29 0 548.55 0.26 ;
        END
    END A_BM[43]
    PIN A_BM[20]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  235.93 0 236.19 0.26 ;
        END
    END A_BM[20]
    PIN A_BIST_BM[43]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  549.665 0 549.925 0.26 ;
        END
    END A_BIST_BM[43]
    PIN A_BIST_BM[20]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  234.555 0 234.815 0.26 ;
        END
    END A_BIST_BM[20]
    PIN A_DOUT[43]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  548.8 0 549.06 0.26 ;
        END
    END A_DOUT[43]
    PIN A_DOUT[20]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  235.42 0 235.68 0.26 ;
        END
    END A_DOUT[20]
    PIN A_DIN[44]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  567.37 0 567.63 0.26 ;
        END
    END A_DIN[44]
    PIN A_DIN[19]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  216.85 0 217.11 0.26 ;
        END
    END A_DIN[19]
    PIN A_BIST_DIN[44]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  566.515 0 566.775 0.26 ;
        END
    END A_BIST_DIN[44]
    PIN A_BIST_DIN[19]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  217.705 0 217.965 0.26 ;
        END
    END A_BIST_DIN[19]
    PIN A_BM[44]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  559.53 0 559.79 0.26 ;
        END
    END A_BM[44]
    PIN A_BM[19]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  224.69 0 224.95 0.26 ;
        END
    END A_BM[19]
    PIN A_BIST_BM[44]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  560.905 0 561.165 0.26 ;
        END
    END A_BIST_BM[44]
    PIN A_BIST_BM[19]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  223.315 0 223.575 0.26 ;
        END
    END A_BIST_BM[19]
    PIN A_DOUT[44]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  560.04 0 560.3 0.26 ;
        END
    END A_DOUT[44]
    PIN A_DOUT[19]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  224.18 0 224.44 0.26 ;
        END
    END A_DOUT[19]
    PIN A_DIN[45]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  578.61 0 578.87 0.26 ;
        END
    END A_DIN[45]
    PIN A_DIN[18]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  205.61 0 205.87 0.26 ;
        END
    END A_DIN[18]
    PIN A_BIST_DIN[45]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  577.755 0 578.015 0.26 ;
        END
    END A_BIST_DIN[45]
    PIN A_BIST_DIN[18]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  206.465 0 206.725 0.26 ;
        END
    END A_BIST_DIN[18]
    PIN A_BM[45]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  570.77 0 571.03 0.26 ;
        END
    END A_BM[45]
    PIN A_BM[18]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  213.45 0 213.71 0.26 ;
        END
    END A_BM[18]
    PIN A_BIST_BM[45]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  572.145 0 572.405 0.26 ;
        END
    END A_BIST_BM[45]
    PIN A_BIST_BM[18]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  212.075 0 212.335 0.26 ;
        END
    END A_BIST_BM[18]
    PIN A_DOUT[45]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  571.28 0 571.54 0.26 ;
        END
    END A_DOUT[45]
    PIN A_DOUT[18]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  212.94 0 213.2 0.26 ;
        END
    END A_DOUT[18]
    PIN A_DIN[46]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  589.85 0 590.11 0.26 ;
        END
    END A_DIN[46]
    PIN A_DIN[17]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  194.37 0 194.63 0.26 ;
        END
    END A_DIN[17]
    PIN A_BIST_DIN[46]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  588.995 0 589.255 0.26 ;
        END
    END A_BIST_DIN[46]
    PIN A_BIST_DIN[17]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  195.225 0 195.485 0.26 ;
        END
    END A_BIST_DIN[17]
    PIN A_BM[46]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  582.01 0 582.27 0.26 ;
        END
    END A_BM[46]
    PIN A_BM[17]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  202.21 0 202.47 0.26 ;
        END
    END A_BM[17]
    PIN A_BIST_BM[46]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  583.385 0 583.645 0.26 ;
        END
    END A_BIST_BM[46]
    PIN A_BIST_BM[17]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  200.835 0 201.095 0.26 ;
        END
    END A_BIST_BM[17]
    PIN A_DOUT[46]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  582.52 0 582.78 0.26 ;
        END
    END A_DOUT[46]
    PIN A_DOUT[17]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  201.7 0 201.96 0.26 ;
        END
    END A_DOUT[17]
    PIN A_DIN[47]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  601.09 0 601.35 0.26 ;
        END
    END A_DIN[47]
    PIN A_DIN[16]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  183.13 0 183.39 0.26 ;
        END
    END A_DIN[16]
    PIN A_BIST_DIN[47]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  600.235 0 600.495 0.26 ;
        END
    END A_BIST_DIN[47]
    PIN A_BIST_DIN[16]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  183.985 0 184.245 0.26 ;
        END
    END A_BIST_DIN[16]
    PIN A_BM[47]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  593.25 0 593.51 0.26 ;
        END
    END A_BM[47]
    PIN A_BM[16]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  190.97 0 191.23 0.26 ;
        END
    END A_BM[16]
    PIN A_BIST_BM[47]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  594.625 0 594.885 0.26 ;
        END
    END A_BIST_BM[47]
    PIN A_BIST_BM[16]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  189.595 0 189.855 0.26 ;
        END
    END A_BIST_BM[16]
    PIN A_DOUT[47]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  593.76 0 594.02 0.26 ;
        END
    END A_DOUT[47]
    PIN A_DOUT[16]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  190.46 0 190.72 0.26 ;
        END
    END A_DOUT[16]
    PIN A_DIN[48]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  612.33 0 612.59 0.26 ;
        END
    END A_DIN[48]
    PIN A_DIN[15]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  171.89 0 172.15 0.26 ;
        END
    END A_DIN[15]
    PIN A_BIST_DIN[48]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  611.475 0 611.735 0.26 ;
        END
    END A_BIST_DIN[48]
    PIN A_BIST_DIN[15]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  172.745 0 173.005 0.26 ;
        END
    END A_BIST_DIN[15]
    PIN A_BM[48]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  604.49 0 604.75 0.26 ;
        END
    END A_BM[48]
    PIN A_BM[15]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  179.73 0 179.99 0.26 ;
        END
    END A_BM[15]
    PIN A_BIST_BM[48]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  605.865 0 606.125 0.26 ;
        END
    END A_BIST_BM[48]
    PIN A_BIST_BM[15]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  178.355 0 178.615 0.26 ;
        END
    END A_BIST_BM[15]
    PIN A_DOUT[48]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  605 0 605.26 0.26 ;
        END
    END A_DOUT[48]
    PIN A_DOUT[15]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  179.22 0 179.48 0.26 ;
        END
    END A_DOUT[15]
    PIN A_DIN[49]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  623.57 0 623.83 0.26 ;
        END
    END A_DIN[49]
    PIN A_DIN[14]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  160.65 0 160.91 0.26 ;
        END
    END A_DIN[14]
    PIN A_BIST_DIN[49]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  622.715 0 622.975 0.26 ;
        END
    END A_BIST_DIN[49]
    PIN A_BIST_DIN[14]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  161.505 0 161.765 0.26 ;
        END
    END A_BIST_DIN[14]
    PIN A_BM[49]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  615.73 0 615.99 0.26 ;
        END
    END A_BM[49]
    PIN A_BM[14]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  168.49 0 168.75 0.26 ;
        END
    END A_BM[14]
    PIN A_BIST_BM[49]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  617.105 0 617.365 0.26 ;
        END
    END A_BIST_BM[49]
    PIN A_BIST_BM[14]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  167.115 0 167.375 0.26 ;
        END
    END A_BIST_BM[14]
    PIN A_DOUT[49]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  616.24 0 616.5 0.26 ;
        END
    END A_DOUT[49]
    PIN A_DOUT[14]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  167.98 0 168.24 0.26 ;
        END
    END A_DOUT[14]
    PIN A_DIN[50]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  634.81 0 635.07 0.26 ;
        END
    END A_DIN[50]
    PIN A_DIN[13]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  149.41 0 149.67 0.26 ;
        END
    END A_DIN[13]
    PIN A_BIST_DIN[50]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  633.955 0 634.215 0.26 ;
        END
    END A_BIST_DIN[50]
    PIN A_BIST_DIN[13]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  150.265 0 150.525 0.26 ;
        END
    END A_BIST_DIN[13]
    PIN A_BM[50]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  626.97 0 627.23 0.26 ;
        END
    END A_BM[50]
    PIN A_BM[13]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  157.25 0 157.51 0.26 ;
        END
    END A_BM[13]
    PIN A_BIST_BM[50]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  628.345 0 628.605 0.26 ;
        END
    END A_BIST_BM[50]
    PIN A_BIST_BM[13]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  155.875 0 156.135 0.26 ;
        END
    END A_BIST_BM[13]
    PIN A_DOUT[50]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  627.48 0 627.74 0.26 ;
        END
    END A_DOUT[50]
    PIN A_DOUT[13]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  156.74 0 157 0.26 ;
        END
    END A_DOUT[13]
    PIN A_DIN[51]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  646.05 0 646.31 0.26 ;
        END
    END A_DIN[51]
    PIN A_DIN[12]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  138.17 0 138.43 0.26 ;
        END
    END A_DIN[12]
    PIN A_BIST_DIN[51]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  645.195 0 645.455 0.26 ;
        END
    END A_BIST_DIN[51]
    PIN A_BIST_DIN[12]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  139.025 0 139.285 0.26 ;
        END
    END A_BIST_DIN[12]
    PIN A_BM[51]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  638.21 0 638.47 0.26 ;
        END
    END A_BM[51]
    PIN A_BM[12]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  146.01 0 146.27 0.26 ;
        END
    END A_BM[12]
    PIN A_BIST_BM[51]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  639.585 0 639.845 0.26 ;
        END
    END A_BIST_BM[51]
    PIN A_BIST_BM[12]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  144.635 0 144.895 0.26 ;
        END
    END A_BIST_BM[12]
    PIN A_DOUT[51]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  638.72 0 638.98 0.26 ;
        END
    END A_DOUT[51]
    PIN A_DOUT[12]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  145.5 0 145.76 0.26 ;
        END
    END A_DOUT[12]
    PIN A_DIN[52]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  657.29 0 657.55 0.26 ;
        END
    END A_DIN[52]
    PIN A_DIN[11]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  126.93 0 127.19 0.26 ;
        END
    END A_DIN[11]
    PIN A_BIST_DIN[52]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  656.435 0 656.695 0.26 ;
        END
    END A_BIST_DIN[52]
    PIN A_BIST_DIN[11]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  127.785 0 128.045 0.26 ;
        END
    END A_BIST_DIN[11]
    PIN A_BM[52]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  649.45 0 649.71 0.26 ;
        END
    END A_BM[52]
    PIN A_BM[11]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  134.77 0 135.03 0.26 ;
        END
    END A_BM[11]
    PIN A_BIST_BM[52]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  650.825 0 651.085 0.26 ;
        END
    END A_BIST_BM[52]
    PIN A_BIST_BM[11]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  133.395 0 133.655 0.26 ;
        END
    END A_BIST_BM[11]
    PIN A_DOUT[52]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  649.96 0 650.22 0.26 ;
        END
    END A_DOUT[52]
    PIN A_DOUT[11]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  134.26 0 134.52 0.26 ;
        END
    END A_DOUT[11]
    PIN A_DIN[53]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  668.53 0 668.79 0.26 ;
        END
    END A_DIN[53]
    PIN A_DIN[10]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  115.69 0 115.95 0.26 ;
        END
    END A_DIN[10]
    PIN A_BIST_DIN[53]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  667.675 0 667.935 0.26 ;
        END
    END A_BIST_DIN[53]
    PIN A_BIST_DIN[10]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  116.545 0 116.805 0.26 ;
        END
    END A_BIST_DIN[10]
    PIN A_BM[53]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  660.69 0 660.95 0.26 ;
        END
    END A_BM[53]
    PIN A_BM[10]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  123.53 0 123.79 0.26 ;
        END
    END A_BM[10]
    PIN A_BIST_BM[53]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  662.065 0 662.325 0.26 ;
        END
    END A_BIST_BM[53]
    PIN A_BIST_BM[10]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  122.155 0 122.415 0.26 ;
        END
    END A_BIST_BM[10]
    PIN A_DOUT[53]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  661.2 0 661.46 0.26 ;
        END
    END A_DOUT[53]
    PIN A_DOUT[10]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  123.02 0 123.28 0.26 ;
        END
    END A_DOUT[10]
    PIN A_DIN[54]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  679.77 0 680.03 0.26 ;
        END
    END A_DIN[54]
    PIN A_DIN[9]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  104.45 0 104.71 0.26 ;
        END
    END A_DIN[9]
    PIN A_BIST_DIN[54]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  678.915 0 679.175 0.26 ;
        END
    END A_BIST_DIN[54]
    PIN A_BIST_DIN[9]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  105.305 0 105.565 0.26 ;
        END
    END A_BIST_DIN[9]
    PIN A_BM[54]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  671.93 0 672.19 0.26 ;
        END
    END A_BM[54]
    PIN A_BM[9]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  112.29 0 112.55 0.26 ;
        END
    END A_BM[9]
    PIN A_BIST_BM[54]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  673.305 0 673.565 0.26 ;
        END
    END A_BIST_BM[54]
    PIN A_BIST_BM[9]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  110.915 0 111.175 0.26 ;
        END
    END A_BIST_BM[9]
    PIN A_DOUT[54]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  672.44 0 672.7 0.26 ;
        END
    END A_DOUT[54]
    PIN A_DOUT[9]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  111.78 0 112.04 0.26 ;
        END
    END A_DOUT[9]
    PIN A_DIN[55]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  691.01 0 691.27 0.26 ;
        END
    END A_DIN[55]
    PIN A_DIN[8]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  93.21 0 93.47 0.26 ;
        END
    END A_DIN[8]
    PIN A_BIST_DIN[55]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  690.155 0 690.415 0.26 ;
        END
    END A_BIST_DIN[55]
    PIN A_BIST_DIN[8]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  94.065 0 94.325 0.26 ;
        END
    END A_BIST_DIN[8]
    PIN A_BM[55]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  683.17 0 683.43 0.26 ;
        END
    END A_BM[55]
    PIN A_BM[8]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  101.05 0 101.31 0.26 ;
        END
    END A_BM[8]
    PIN A_BIST_BM[55]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  684.545 0 684.805 0.26 ;
        END
    END A_BIST_BM[55]
    PIN A_BIST_BM[8]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  99.675 0 99.935 0.26 ;
        END
    END A_BIST_BM[8]
    PIN A_DOUT[55]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  683.68 0 683.94 0.26 ;
        END
    END A_DOUT[55]
    PIN A_DOUT[8]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  100.54 0 100.8 0.26 ;
        END
    END A_DOUT[8]
    PIN A_DIN[56]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  702.25 0 702.51 0.26 ;
        END
    END A_DIN[56]
    PIN A_DIN[7]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  81.97 0 82.23 0.26 ;
        END
    END A_DIN[7]
    PIN A_BIST_DIN[56]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  701.395 0 701.655 0.26 ;
        END
    END A_BIST_DIN[56]
    PIN A_BIST_DIN[7]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  82.825 0 83.085 0.26 ;
        END
    END A_BIST_DIN[7]
    PIN A_BM[56]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  694.41 0 694.67 0.26 ;
        END
    END A_BM[56]
    PIN A_BM[7]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  89.81 0 90.07 0.26 ;
        END
    END A_BM[7]
    PIN A_BIST_BM[56]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  695.785 0 696.045 0.26 ;
        END
    END A_BIST_BM[56]
    PIN A_BIST_BM[7]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  88.435 0 88.695 0.26 ;
        END
    END A_BIST_BM[7]
    PIN A_DOUT[56]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  694.92 0 695.18 0.26 ;
        END
    END A_DOUT[56]
    PIN A_DOUT[7]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  89.3 0 89.56 0.26 ;
        END
    END A_DOUT[7]
    PIN A_DIN[57]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  713.49 0 713.75 0.26 ;
        END
    END A_DIN[57]
    PIN A_DIN[6]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  70.73 0 70.99 0.26 ;
        END
    END A_DIN[6]
    PIN A_BIST_DIN[57]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  712.635 0 712.895 0.26 ;
        END
    END A_BIST_DIN[57]
    PIN A_BIST_DIN[6]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  71.585 0 71.845 0.26 ;
        END
    END A_BIST_DIN[6]
    PIN A_BM[57]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  705.65 0 705.91 0.26 ;
        END
    END A_BM[57]
    PIN A_BM[6]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  78.57 0 78.83 0.26 ;
        END
    END A_BM[6]
    PIN A_BIST_BM[57]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  707.025 0 707.285 0.26 ;
        END
    END A_BIST_BM[57]
    PIN A_BIST_BM[6]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  77.195 0 77.455 0.26 ;
        END
    END A_BIST_BM[6]
    PIN A_DOUT[57]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  706.16 0 706.42 0.26 ;
        END
    END A_DOUT[57]
    PIN A_DOUT[6]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  78.06 0 78.32 0.26 ;
        END
    END A_DOUT[6]
    PIN A_DIN[58]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  724.73 0 724.99 0.26 ;
        END
    END A_DIN[58]
    PIN A_DIN[5]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  59.49 0 59.75 0.26 ;
        END
    END A_DIN[5]
    PIN A_BIST_DIN[58]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  723.875 0 724.135 0.26 ;
        END
    END A_BIST_DIN[58]
    PIN A_BIST_DIN[5]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  60.345 0 60.605 0.26 ;
        END
    END A_BIST_DIN[5]
    PIN A_BM[58]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  716.89 0 717.15 0.26 ;
        END
    END A_BM[58]
    PIN A_BM[5]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  67.33 0 67.59 0.26 ;
        END
    END A_BM[5]
    PIN A_BIST_BM[58]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  718.265 0 718.525 0.26 ;
        END
    END A_BIST_BM[58]
    PIN A_BIST_BM[5]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  65.955 0 66.215 0.26 ;
        END
    END A_BIST_BM[5]
    PIN A_DOUT[58]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  717.4 0 717.66 0.26 ;
        END
    END A_DOUT[58]
    PIN A_DOUT[5]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  66.82 0 67.08 0.26 ;
        END
    END A_DOUT[5]
    PIN A_DIN[59]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  735.97 0 736.23 0.26 ;
        END
    END A_DIN[59]
    PIN A_DIN[4]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  48.25 0 48.51 0.26 ;
        END
    END A_DIN[4]
    PIN A_BIST_DIN[59]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  735.115 0 735.375 0.26 ;
        END
    END A_BIST_DIN[59]
    PIN A_BIST_DIN[4]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  49.105 0 49.365 0.26 ;
        END
    END A_BIST_DIN[4]
    PIN A_BM[59]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  728.13 0 728.39 0.26 ;
        END
    END A_BM[59]
    PIN A_BM[4]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  56.09 0 56.35 0.26 ;
        END
    END A_BM[4]
    PIN A_BIST_BM[59]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  729.505 0 729.765 0.26 ;
        END
    END A_BIST_BM[59]
    PIN A_BIST_BM[4]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  54.715 0 54.975 0.26 ;
        END
    END A_BIST_BM[4]
    PIN A_DOUT[59]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  728.64 0 728.9 0.26 ;
        END
    END A_DOUT[59]
    PIN A_DOUT[4]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  55.58 0 55.84 0.26 ;
        END
    END A_DOUT[4]
    PIN A_DIN[60]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  747.21 0 747.47 0.26 ;
        END
    END A_DIN[60]
    PIN A_DIN[3]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  37.01 0 37.27 0.26 ;
        END
    END A_DIN[3]
    PIN A_BIST_DIN[60]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  746.355 0 746.615 0.26 ;
        END
    END A_BIST_DIN[60]
    PIN A_BIST_DIN[3]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  37.865 0 38.125 0.26 ;
        END
    END A_BIST_DIN[3]
    PIN A_BM[60]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  739.37 0 739.63 0.26 ;
        END
    END A_BM[60]
    PIN A_BM[3]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  44.85 0 45.11 0.26 ;
        END
    END A_BM[3]
    PIN A_BIST_BM[60]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  740.745 0 741.005 0.26 ;
        END
    END A_BIST_BM[60]
    PIN A_BIST_BM[3]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  43.475 0 43.735 0.26 ;
        END
    END A_BIST_BM[3]
    PIN A_DOUT[60]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  739.88 0 740.14 0.26 ;
        END
    END A_DOUT[60]
    PIN A_DOUT[3]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  44.34 0 44.6 0.26 ;
        END
    END A_DOUT[3]
    PIN A_DIN[61]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  758.45 0 758.71 0.26 ;
        END
    END A_DIN[61]
    PIN A_DIN[2]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  25.77 0 26.03 0.26 ;
        END
    END A_DIN[2]
    PIN A_BIST_DIN[61]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  757.595 0 757.855 0.26 ;
        END
    END A_BIST_DIN[61]
    PIN A_BIST_DIN[2]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  26.625 0 26.885 0.26 ;
        END
    END A_BIST_DIN[2]
    PIN A_BM[61]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  750.61 0 750.87 0.26 ;
        END
    END A_BM[61]
    PIN A_BM[2]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  33.61 0 33.87 0.26 ;
        END
    END A_BM[2]
    PIN A_BIST_BM[61]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  751.985 0 752.245 0.26 ;
        END
    END A_BIST_BM[61]
    PIN A_BIST_BM[2]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  32.235 0 32.495 0.26 ;
        END
    END A_BIST_BM[2]
    PIN A_DOUT[61]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  751.12 0 751.38 0.26 ;
        END
    END A_DOUT[61]
    PIN A_DOUT[2]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  33.1 0 33.36 0.26 ;
        END
    END A_DOUT[2]
    PIN A_DIN[62]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  769.69 0 769.95 0.26 ;
        END
    END A_DIN[62]
    PIN A_DIN[1]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  14.53 0 14.79 0.26 ;
        END
    END A_DIN[1]
    PIN A_BIST_DIN[62]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  768.835 0 769.095 0.26 ;
        END
    END A_BIST_DIN[62]
    PIN A_BIST_DIN[1]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  15.385 0 15.645 0.26 ;
        END
    END A_BIST_DIN[1]
    PIN A_BM[62]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  761.85 0 762.11 0.26 ;
        END
    END A_BM[62]
    PIN A_BM[1]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  22.37 0 22.63 0.26 ;
        END
    END A_BM[1]
    PIN A_BIST_BM[62]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  763.225 0 763.485 0.26 ;
        END
    END A_BIST_BM[62]
    PIN A_BIST_BM[1]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  20.995 0 21.255 0.26 ;
        END
    END A_BIST_BM[1]
    PIN A_DOUT[62]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  762.36 0 762.62 0.26 ;
        END
    END A_DOUT[62]
    PIN A_DOUT[1]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  21.86 0 22.12 0.26 ;
        END
    END A_DOUT[1]
    PIN A_DIN[63]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  780.93 0 781.19 0.26 ;
        END
    END A_DIN[63]
    PIN A_DIN[0]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.83819 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  3.29 0 3.55 0.26 ;
        END
    END A_DIN[0]
    PIN A_BIST_DIN[63]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  780.075 0 780.335 0.26 ;
        END
    END A_BIST_DIN[63]
    PIN A_BIST_DIN[0]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 9.36594 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  4.145 0 4.405 0.26 ;
        END
    END A_BIST_DIN[0]
    PIN A_BM[63]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  773.09 0 773.35 0.26 ;
        END
    END A_BM[63]
    PIN A_BM[0]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 4.49838 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  11.13 0 11.39 0.26 ;
        END
    END A_BM[0]
    PIN A_BIST_BM[63]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  774.465 0 774.725 0.26 ;
        END
    END A_BIST_BM[63]
    PIN A_BIST_BM[0]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 5.05527 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  9.755 0 10.015 0.26 ;
        END
    END A_BIST_BM[0]
    PIN A_DOUT[63]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  773.6 0 773.86 0.26 ;
        END
    END A_DOUT[63]
    PIN A_DOUT[0]
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
        ANTENNADIFFAREA 0.988 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  10.62 0 10.88 0.26 ;
        END
    END A_DOUT[0]
    PIN A_ADDR[0]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 8.9011 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 45.2233 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  388.44 0 388.7 0.26 ;
        END
    END A_ADDR[0]
    PIN A_BIST_ADDR[0]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 9.6967 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 49.1845 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  393.03 0 393.29 0.26 ;
        END
    END A_BIST_ADDR[0]
    PIN A_ADDR[1]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 7.774 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 39.657 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  387.93 0 388.19 0.26 ;
        END
    END A_ADDR[1]
    PIN A_BIST_ADDR[1]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 8.5696 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 43.6181 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  392.52 0 392.78 0.26 ;
        END
    END A_BIST_ADDR[1]
    PIN A_ADDR[2]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 10.6327 LAYER Metal2 ;
        ANTENNAPARTIALMETALAREA 1.5246 LAYER Metal3 ;
        ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
        ANTENNAMAXAREACAR 9.41598 LAYER Metal3 ;
        PORT
            LAYER Metal2 ;
              RECT  396.09 0 396.35 0.26 ;
        END
    END A_ADDR[2]
    PIN A_BIST_ADDR[2]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 10.6327 LAYER Metal2 ;
        ANTENNAPARTIALMETALAREA 1.0962 LAYER Metal3 ;
        ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
        ANTENNAMAXAREACAR 7.81379 LAYER Metal3 ;
        PORT
            LAYER Metal2 ;
              RECT  396.6 0 396.86 0.26 ;
        END
    END A_BIST_ADDR[2]
    PIN A_ADDR[3]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 10.6327 LAYER Metal2 ;
        ANTENNAPARTIALMETALAREA 3.8367 LAYER Metal3 ;
        ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
        ANTENNAMAXAREACAR 20.9276 LAYER Metal3 ;
        PORT
            LAYER Metal2 ;
              RECT  395.07 0 395.33 0.26 ;
        END
    END A_ADDR[3]
    PIN A_BIST_ADDR[3]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 10.6327 LAYER Metal2 ;
        ANTENNAPARTIALMETALAREA 3.5175 LAYER Metal3 ;
        ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
        ANTENNAMAXAREACAR 19.8691 LAYER Metal3 ;
        PORT
            LAYER Metal2 ;
              RECT  395.58 0 395.84 0.26 ;
        END
    END A_BIST_ADDR[3]
    PIN A_ADDR[4]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 12.1979 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 61.6375 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  398.64 0 398.9 0.26 ;
        END
    END A_ADDR[4]
    PIN A_BIST_ADDR[4]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 11.9327 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 60.3172 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  398.13 0 398.39 0.26 ;
        END
    END A_BIST_ADDR[4]
    PIN A_ADDR[5]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 13.9269 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 70.246 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  397.62 0 397.88 0.26 ;
        END
    END A_ADDR[5]
    PIN A_BIST_ADDR[5]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 13.6617 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 68.9256 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  397.11 0 397.37 0.26 ;
        END
    END A_BIST_ADDR[5]
    PIN A_ADDR[6]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 10.9525 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 55.4369 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  376.2 0 376.46 0.26 ;
        END
    END A_ADDR[6]
    PIN A_BIST_ADDR[6]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 10.6771 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 54.0657 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  376.71 0 376.97 0.26 ;
        END
    END A_BIST_ADDR[6]
    PIN A_ADDR[7]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 12.4163 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 62.7249 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  377.22 0 377.48 0.26 ;
        END
    END A_ADDR[7]
    PIN A_BIST_ADDR[7]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 12.1511 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 61.4045 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  377.73 0 377.99 0.26 ;
        END
    END A_BIST_ADDR[7]
    PIN A_ADDR[8]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 10.3675 LAYER Metal2 ;
        ANTENNAPARTIALMETALAREA 1.5897 LAYER Metal3 ;
        ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
        ANTENNAMAXAREACAR 9.7401 LAYER Metal3 ;
        PORT
            LAYER Metal2 ;
              RECT  406.29 0 406.55 0.26 ;
        END
    END A_ADDR[8]
    PIN A_BIST_ADDR[8]
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 10.3675 LAYER Metal2 ;
        ANTENNAPARTIALMETALAREA 1.3755 LAYER Metal3 ;
        ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
        ANTENNAMAXAREACAR 9.20438 LAYER Metal3 ;
        PORT
            LAYER Metal2 ;
              RECT  406.8 0 407.06 0.26 ;
        END
    END A_BIST_ADDR[8]
    PIN A_CLK
        DIRECTION INPUT ; 
        USE CLOCK ; 
        ANTENNAPARTIALMETALAREA 4.0547 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 21.0939 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  386.4 0 386.66 0.26 ;
        END
    END A_CLK
    PIN A_REN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.99505 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 20.7969 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  389.97 0 390.23 0.26 ;
        END
    END A_REN
    PIN A_WEN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 15.2686 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  389.46 0 389.72 0.26 ;
        END
    END A_WEN
    PIN A_MEN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.0247 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 15.9656 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  386.91 0 387.17 0.26 ;
        END
    END A_MEN
    PIN A_DLY
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 6.058 LAYER Metal2 ;
        ANTENNAGATEAREA 0.3367 LAYER Metal2 ;
        ANTENNAMAXAREACAR 18.5328 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  408.33 0 408.59 0.26 ;
        END
    END A_DLY
    PIN A_BIST_EN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 3.9871 LAYER Metal2 ;
        ANTENNAPARTIALMETALAREA 382.413 LAYER Metal3 ;
        ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
        ANTENNAGATEAREA 1.43 LAYER Metal2 ;
        ANTENNAGATEAREA 50.4075 LAYER Metal3 ;
        ANTENNAMAXAREACAR 3.21364 LAYER Metal2 ;
        ANTENNAMAXAREACAR 17.8592 LAYER Metal3 ;
        ANTENNAMAXCUTCAR 0.151469 LAYER Via2 ;
        PORT
            LAYER Metal2 ;
              RECT  388.95 0 389.21 0.26 ;
        END
    END A_BIST_EN
    PIN A_BIST_CLK
        DIRECTION INPUT ; 
        USE CLOCK ; 
        ANTENNAPARTIALMETALAREA 4.1639 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 21.9534 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  384.87 0 385.13 0.26 ;
        END
    END A_BIST_CLK
    PIN A_BIST_REN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 4.1119 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 21.6945 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  391.5 0 391.76 0.26 ;
        END
    END A_BIST_REN
    PIN A_BIST_WEN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 2.9051 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 15.6861 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  390.99 0 391.25 0.26 ;
        END
    END A_BIST_WEN
    PIN A_BIST_MEN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        ANTENNAPARTIALMETALAREA 2.8977 LAYER Metal2 ;
        ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
        ANTENNAMAXAREACAR 15.6492 LAYER Metal2 ;
        PORT
            LAYER Metal2 ;
              RECT  385.38 0 385.64 0.26 ;
        END
    END A_BIST_MEN
    OBS
      LAYER Metal1 ;
        RECT  0 0 784.48 191.34 ;
      LAYER Metal2 ;
        RECT  0.105 45.465 0.305 191.315 ;
        RECT  1.1 190.585 1.3 191.315 ;
        RECT  3.29 0.52 3.55 5.16 ;
        RECT  2.77 4.9 3.55 5.16 ;
        RECT  2.77 4.9 3.03 6.64 ;
        RECT  1.92 190.585 2.12 191.315 ;
        RECT  2.415 190.585 2.615 191.315 ;
        RECT  2.915 190.585 3.115 191.315 ;
        RECT  3.415 190.585 3.615 191.315 ;
        RECT  3.91 190.585 4.11 191.315 ;
        RECT  4.655 0.17 5.425 0.94 ;
        RECT  4.655 0.17 4.915 12.9 ;
        RECT  5.165 0.17 5.425 12.9 ;
        RECT  4.145 0.52 4.405 5.815 ;
        RECT  4.73 190.585 4.93 191.315 ;
        RECT  5.675 0.17 6.445 0.43 ;
        RECT  5.675 0.17 5.935 11.5 ;
        RECT  6.185 0.17 6.445 11.5 ;
        RECT  5.225 190.585 5.425 191.315 ;
        RECT  5.725 190.585 5.925 191.315 ;
        RECT  6.225 190.585 6.425 191.315 ;
        RECT  7.715 0.17 8.485 0.43 ;
        RECT  7.715 0.17 7.975 10.48 ;
        RECT  8.225 0.17 8.485 10.99 ;
        RECT  6.72 190.585 6.92 191.315 ;
        RECT  7.54 190.585 7.74 191.315 ;
        RECT  8.735 0.17 9.505 0.94 ;
        RECT  8.735 0.17 8.995 8.7 ;
        RECT  9.245 0.17 9.505 12.9 ;
        RECT  8.035 190.585 8.235 191.315 ;
        RECT  8.535 190.585 8.735 191.315 ;
        RECT  9.035 190.585 9.235 191.315 ;
        RECT  9.53 190.585 9.73 191.315 ;
        RECT  9.755 0.52 10.015 2.485 ;
        RECT  10.35 190.585 10.55 191.315 ;
        RECT  10.62 0.52 10.88 14.11 ;
        RECT  10.845 190.585 11.045 191.315 ;
        RECT  11.13 0.52 11.39 2.335 ;
        RECT  11.345 190.585 11.545 191.315 ;
        RECT  11.845 190.585 12.045 191.315 ;
        RECT  12.34 190.585 12.54 191.315 ;
        RECT  14.53 0.52 14.79 5.16 ;
        RECT  14.01 4.9 14.79 5.16 ;
        RECT  14.01 4.9 14.27 6.64 ;
        RECT  13.16 190.585 13.36 191.315 ;
        RECT  13.655 190.585 13.855 191.315 ;
        RECT  14.155 190.585 14.355 191.315 ;
        RECT  14.655 190.585 14.855 191.315 ;
        RECT  15.15 190.585 15.35 191.315 ;
        RECT  15.895 0.17 16.665 0.94 ;
        RECT  15.895 0.17 16.155 12.9 ;
        RECT  16.405 0.17 16.665 12.9 ;
        RECT  15.385 0.52 15.645 5.815 ;
        RECT  15.97 190.585 16.17 191.315 ;
        RECT  16.915 0.17 17.685 0.43 ;
        RECT  16.915 0.17 17.175 11.5 ;
        RECT  17.425 0.17 17.685 11.5 ;
        RECT  16.465 190.585 16.665 191.315 ;
        RECT  16.965 190.585 17.165 191.315 ;
        RECT  17.465 190.585 17.665 191.315 ;
        RECT  18.955 0.17 19.725 0.43 ;
        RECT  18.955 0.17 19.215 10.48 ;
        RECT  19.465 0.17 19.725 10.99 ;
        RECT  17.96 190.585 18.16 191.315 ;
        RECT  18.78 190.585 18.98 191.315 ;
        RECT  19.975 0.17 20.745 0.94 ;
        RECT  19.975 0.17 20.235 8.7 ;
        RECT  20.485 0.17 20.745 12.9 ;
        RECT  19.275 190.585 19.475 191.315 ;
        RECT  19.775 190.585 19.975 191.315 ;
        RECT  20.275 190.585 20.475 191.315 ;
        RECT  20.77 190.585 20.97 191.315 ;
        RECT  20.995 0.52 21.255 2.485 ;
        RECT  21.59 190.585 21.79 191.315 ;
        RECT  21.86 0.52 22.12 14.11 ;
        RECT  22.085 190.585 22.285 191.315 ;
        RECT  22.37 0.52 22.63 2.335 ;
        RECT  22.585 190.585 22.785 191.315 ;
        RECT  23.085 190.585 23.285 191.315 ;
        RECT  23.58 190.585 23.78 191.315 ;
        RECT  25.77 0.52 26.03 5.16 ;
        RECT  25.25 4.9 26.03 5.16 ;
        RECT  25.25 4.9 25.51 6.64 ;
        RECT  24.4 190.585 24.6 191.315 ;
        RECT  24.895 190.585 25.095 191.315 ;
        RECT  25.395 190.585 25.595 191.315 ;
        RECT  25.895 190.585 26.095 191.315 ;
        RECT  26.39 190.585 26.59 191.315 ;
        RECT  27.135 0.17 27.905 0.94 ;
        RECT  27.135 0.17 27.395 12.9 ;
        RECT  27.645 0.17 27.905 12.9 ;
        RECT  26.625 0.52 26.885 5.815 ;
        RECT  27.21 190.585 27.41 191.315 ;
        RECT  28.155 0.17 28.925 0.43 ;
        RECT  28.155 0.17 28.415 11.5 ;
        RECT  28.665 0.17 28.925 11.5 ;
        RECT  27.705 190.585 27.905 191.315 ;
        RECT  28.205 190.585 28.405 191.315 ;
        RECT  28.705 190.585 28.905 191.315 ;
        RECT  30.195 0.17 30.965 0.43 ;
        RECT  30.195 0.17 30.455 10.48 ;
        RECT  30.705 0.17 30.965 10.99 ;
        RECT  29.2 190.585 29.4 191.315 ;
        RECT  30.02 190.585 30.22 191.315 ;
        RECT  31.215 0.17 31.985 0.94 ;
        RECT  31.215 0.17 31.475 8.7 ;
        RECT  31.725 0.17 31.985 12.9 ;
        RECT  30.515 190.585 30.715 191.315 ;
        RECT  31.015 190.585 31.215 191.315 ;
        RECT  31.515 190.585 31.715 191.315 ;
        RECT  32.01 190.585 32.21 191.315 ;
        RECT  32.235 0.52 32.495 2.485 ;
        RECT  32.83 190.585 33.03 191.315 ;
        RECT  33.1 0.52 33.36 14.11 ;
        RECT  33.325 190.585 33.525 191.315 ;
        RECT  33.61 0.52 33.87 2.335 ;
        RECT  33.825 190.585 34.025 191.315 ;
        RECT  34.325 190.585 34.525 191.315 ;
        RECT  34.82 190.585 35.02 191.315 ;
        RECT  37.01 0.52 37.27 5.16 ;
        RECT  36.49 4.9 37.27 5.16 ;
        RECT  36.49 4.9 36.75 6.64 ;
        RECT  35.64 190.585 35.84 191.315 ;
        RECT  36.135 190.585 36.335 191.315 ;
        RECT  36.635 190.585 36.835 191.315 ;
        RECT  37.135 190.585 37.335 191.315 ;
        RECT  37.63 190.585 37.83 191.315 ;
        RECT  38.375 0.17 39.145 0.94 ;
        RECT  38.375 0.17 38.635 12.9 ;
        RECT  38.885 0.17 39.145 12.9 ;
        RECT  37.865 0.52 38.125 5.815 ;
        RECT  38.45 190.585 38.65 191.315 ;
        RECT  39.395 0.17 40.165 0.43 ;
        RECT  39.395 0.17 39.655 11.5 ;
        RECT  39.905 0.17 40.165 11.5 ;
        RECT  38.945 190.585 39.145 191.315 ;
        RECT  39.445 190.585 39.645 191.315 ;
        RECT  39.945 190.585 40.145 191.315 ;
        RECT  41.435 0.17 42.205 0.43 ;
        RECT  41.435 0.17 41.695 10.48 ;
        RECT  41.945 0.17 42.205 10.99 ;
        RECT  40.44 190.585 40.64 191.315 ;
        RECT  41.26 190.585 41.46 191.315 ;
        RECT  42.455 0.17 43.225 0.94 ;
        RECT  42.455 0.17 42.715 8.7 ;
        RECT  42.965 0.17 43.225 12.9 ;
        RECT  41.755 190.585 41.955 191.315 ;
        RECT  42.255 190.585 42.455 191.315 ;
        RECT  42.755 190.585 42.955 191.315 ;
        RECT  43.25 190.585 43.45 191.315 ;
        RECT  43.475 0.52 43.735 2.485 ;
        RECT  44.07 190.585 44.27 191.315 ;
        RECT  44.34 0.52 44.6 14.11 ;
        RECT  44.565 190.585 44.765 191.315 ;
        RECT  44.85 0.52 45.11 2.335 ;
        RECT  45.065 190.585 45.265 191.315 ;
        RECT  45.565 190.585 45.765 191.315 ;
        RECT  46.06 190.585 46.26 191.315 ;
        RECT  48.25 0.52 48.51 5.16 ;
        RECT  47.73 4.9 48.51 5.16 ;
        RECT  47.73 4.9 47.99 6.64 ;
        RECT  46.88 190.585 47.08 191.315 ;
        RECT  47.375 190.585 47.575 191.315 ;
        RECT  47.875 190.585 48.075 191.315 ;
        RECT  48.375 190.585 48.575 191.315 ;
        RECT  48.87 190.585 49.07 191.315 ;
        RECT  49.615 0.17 50.385 0.94 ;
        RECT  49.615 0.17 49.875 12.9 ;
        RECT  50.125 0.17 50.385 12.9 ;
        RECT  49.105 0.52 49.365 5.815 ;
        RECT  49.69 190.585 49.89 191.315 ;
        RECT  50.635 0.17 51.405 0.43 ;
        RECT  50.635 0.17 50.895 11.5 ;
        RECT  51.145 0.17 51.405 11.5 ;
        RECT  50.185 190.585 50.385 191.315 ;
        RECT  50.685 190.585 50.885 191.315 ;
        RECT  51.185 190.585 51.385 191.315 ;
        RECT  52.675 0.17 53.445 0.43 ;
        RECT  52.675 0.17 52.935 10.48 ;
        RECT  53.185 0.17 53.445 10.99 ;
        RECT  51.68 190.585 51.88 191.315 ;
        RECT  52.5 190.585 52.7 191.315 ;
        RECT  53.695 0.17 54.465 0.94 ;
        RECT  53.695 0.17 53.955 8.7 ;
        RECT  54.205 0.17 54.465 12.9 ;
        RECT  52.995 190.585 53.195 191.315 ;
        RECT  53.495 190.585 53.695 191.315 ;
        RECT  53.995 190.585 54.195 191.315 ;
        RECT  54.49 190.585 54.69 191.315 ;
        RECT  54.715 0.52 54.975 2.485 ;
        RECT  55.31 190.585 55.51 191.315 ;
        RECT  55.58 0.52 55.84 14.11 ;
        RECT  55.805 190.585 56.005 191.315 ;
        RECT  56.09 0.52 56.35 2.335 ;
        RECT  56.305 190.585 56.505 191.315 ;
        RECT  56.805 190.585 57.005 191.315 ;
        RECT  57.3 190.585 57.5 191.315 ;
        RECT  59.49 0.52 59.75 5.16 ;
        RECT  58.97 4.9 59.75 5.16 ;
        RECT  58.97 4.9 59.23 6.64 ;
        RECT  58.12 190.585 58.32 191.315 ;
        RECT  58.615 190.585 58.815 191.315 ;
        RECT  59.115 190.585 59.315 191.315 ;
        RECT  59.615 190.585 59.815 191.315 ;
        RECT  60.11 190.585 60.31 191.315 ;
        RECT  60.855 0.17 61.625 0.94 ;
        RECT  60.855 0.17 61.115 12.9 ;
        RECT  61.365 0.17 61.625 12.9 ;
        RECT  60.345 0.52 60.605 5.815 ;
        RECT  60.93 190.585 61.13 191.315 ;
        RECT  61.875 0.17 62.645 0.43 ;
        RECT  61.875 0.17 62.135 11.5 ;
        RECT  62.385 0.17 62.645 11.5 ;
        RECT  61.425 190.585 61.625 191.315 ;
        RECT  61.925 190.585 62.125 191.315 ;
        RECT  62.425 190.585 62.625 191.315 ;
        RECT  63.915 0.17 64.685 0.43 ;
        RECT  63.915 0.17 64.175 10.48 ;
        RECT  64.425 0.17 64.685 10.99 ;
        RECT  62.92 190.585 63.12 191.315 ;
        RECT  63.74 190.585 63.94 191.315 ;
        RECT  64.935 0.17 65.705 0.94 ;
        RECT  64.935 0.17 65.195 8.7 ;
        RECT  65.445 0.17 65.705 12.9 ;
        RECT  64.235 190.585 64.435 191.315 ;
        RECT  64.735 190.585 64.935 191.315 ;
        RECT  65.235 190.585 65.435 191.315 ;
        RECT  65.73 190.585 65.93 191.315 ;
        RECT  65.955 0.52 66.215 2.485 ;
        RECT  66.55 190.585 66.75 191.315 ;
        RECT  66.82 0.52 67.08 14.11 ;
        RECT  67.045 190.585 67.245 191.315 ;
        RECT  67.33 0.52 67.59 2.335 ;
        RECT  67.545 190.585 67.745 191.315 ;
        RECT  68.045 190.585 68.245 191.315 ;
        RECT  68.54 190.585 68.74 191.315 ;
        RECT  70.73 0.52 70.99 5.16 ;
        RECT  70.21 4.9 70.99 5.16 ;
        RECT  70.21 4.9 70.47 6.64 ;
        RECT  69.36 190.585 69.56 191.315 ;
        RECT  69.855 190.585 70.055 191.315 ;
        RECT  70.355 190.585 70.555 191.315 ;
        RECT  70.855 190.585 71.055 191.315 ;
        RECT  71.35 190.585 71.55 191.315 ;
        RECT  72.095 0.17 72.865 0.94 ;
        RECT  72.095 0.17 72.355 12.9 ;
        RECT  72.605 0.17 72.865 12.9 ;
        RECT  71.585 0.52 71.845 5.815 ;
        RECT  72.17 190.585 72.37 191.315 ;
        RECT  73.115 0.17 73.885 0.43 ;
        RECT  73.115 0.17 73.375 11.5 ;
        RECT  73.625 0.17 73.885 11.5 ;
        RECT  72.665 190.585 72.865 191.315 ;
        RECT  73.165 190.585 73.365 191.315 ;
        RECT  73.665 190.585 73.865 191.315 ;
        RECT  75.155 0.17 75.925 0.43 ;
        RECT  75.155 0.17 75.415 10.48 ;
        RECT  75.665 0.17 75.925 10.99 ;
        RECT  74.16 190.585 74.36 191.315 ;
        RECT  74.98 190.585 75.18 191.315 ;
        RECT  76.175 0.17 76.945 0.94 ;
        RECT  76.175 0.17 76.435 8.7 ;
        RECT  76.685 0.17 76.945 12.9 ;
        RECT  75.475 190.585 75.675 191.315 ;
        RECT  75.975 190.585 76.175 191.315 ;
        RECT  76.475 190.585 76.675 191.315 ;
        RECT  76.97 190.585 77.17 191.315 ;
        RECT  77.195 0.52 77.455 2.485 ;
        RECT  77.79 190.585 77.99 191.315 ;
        RECT  78.06 0.52 78.32 14.11 ;
        RECT  78.285 190.585 78.485 191.315 ;
        RECT  78.57 0.52 78.83 2.335 ;
        RECT  78.785 190.585 78.985 191.315 ;
        RECT  79.285 190.585 79.485 191.315 ;
        RECT  79.78 190.585 79.98 191.315 ;
        RECT  81.97 0.52 82.23 5.16 ;
        RECT  81.45 4.9 82.23 5.16 ;
        RECT  81.45 4.9 81.71 6.64 ;
        RECT  80.6 190.585 80.8 191.315 ;
        RECT  81.095 190.585 81.295 191.315 ;
        RECT  81.595 190.585 81.795 191.315 ;
        RECT  82.095 190.585 82.295 191.315 ;
        RECT  82.59 190.585 82.79 191.315 ;
        RECT  83.335 0.17 84.105 0.94 ;
        RECT  83.335 0.17 83.595 12.9 ;
        RECT  83.845 0.17 84.105 12.9 ;
        RECT  82.825 0.52 83.085 5.815 ;
        RECT  83.41 190.585 83.61 191.315 ;
        RECT  84.355 0.17 85.125 0.43 ;
        RECT  84.355 0.17 84.615 11.5 ;
        RECT  84.865 0.17 85.125 11.5 ;
        RECT  83.905 190.585 84.105 191.315 ;
        RECT  84.405 190.585 84.605 191.315 ;
        RECT  84.905 190.585 85.105 191.315 ;
        RECT  86.395 0.17 87.165 0.43 ;
        RECT  86.395 0.17 86.655 10.48 ;
        RECT  86.905 0.17 87.165 10.99 ;
        RECT  85.4 190.585 85.6 191.315 ;
        RECT  86.22 190.585 86.42 191.315 ;
        RECT  87.415 0.17 88.185 0.94 ;
        RECT  87.415 0.17 87.675 8.7 ;
        RECT  87.925 0.17 88.185 12.9 ;
        RECT  86.715 190.585 86.915 191.315 ;
        RECT  87.215 190.585 87.415 191.315 ;
        RECT  87.715 190.585 87.915 191.315 ;
        RECT  88.21 190.585 88.41 191.315 ;
        RECT  88.435 0.52 88.695 2.485 ;
        RECT  89.03 190.585 89.23 191.315 ;
        RECT  89.3 0.52 89.56 14.11 ;
        RECT  89.525 190.585 89.725 191.315 ;
        RECT  89.81 0.52 90.07 2.335 ;
        RECT  90.025 190.585 90.225 191.315 ;
        RECT  90.525 190.585 90.725 191.315 ;
        RECT  91.02 190.585 91.22 191.315 ;
        RECT  93.21 0.52 93.47 5.16 ;
        RECT  92.69 4.9 93.47 5.16 ;
        RECT  92.69 4.9 92.95 6.64 ;
        RECT  91.84 190.585 92.04 191.315 ;
        RECT  92.335 190.585 92.535 191.315 ;
        RECT  92.835 190.585 93.035 191.315 ;
        RECT  93.335 190.585 93.535 191.315 ;
        RECT  93.83 190.585 94.03 191.315 ;
        RECT  94.575 0.17 95.345 0.94 ;
        RECT  94.575 0.17 94.835 12.9 ;
        RECT  95.085 0.17 95.345 12.9 ;
        RECT  94.065 0.52 94.325 5.815 ;
        RECT  94.65 190.585 94.85 191.315 ;
        RECT  95.595 0.17 96.365 0.43 ;
        RECT  95.595 0.17 95.855 11.5 ;
        RECT  96.105 0.17 96.365 11.5 ;
        RECT  95.145 190.585 95.345 191.315 ;
        RECT  95.645 190.585 95.845 191.315 ;
        RECT  96.145 190.585 96.345 191.315 ;
        RECT  97.635 0.17 98.405 0.43 ;
        RECT  97.635 0.17 97.895 10.48 ;
        RECT  98.145 0.17 98.405 10.99 ;
        RECT  96.64 190.585 96.84 191.315 ;
        RECT  97.46 190.585 97.66 191.315 ;
        RECT  98.655 0.17 99.425 0.94 ;
        RECT  98.655 0.17 98.915 8.7 ;
        RECT  99.165 0.17 99.425 12.9 ;
        RECT  97.955 190.585 98.155 191.315 ;
        RECT  98.455 190.585 98.655 191.315 ;
        RECT  98.955 190.585 99.155 191.315 ;
        RECT  99.45 190.585 99.65 191.315 ;
        RECT  99.675 0.52 99.935 2.485 ;
        RECT  100.27 190.585 100.47 191.315 ;
        RECT  100.54 0.52 100.8 14.11 ;
        RECT  100.765 190.585 100.965 191.315 ;
        RECT  101.05 0.52 101.31 2.335 ;
        RECT  101.265 190.585 101.465 191.315 ;
        RECT  101.765 190.585 101.965 191.315 ;
        RECT  102.26 190.585 102.46 191.315 ;
        RECT  104.45 0.52 104.71 5.16 ;
        RECT  103.93 4.9 104.71 5.16 ;
        RECT  103.93 4.9 104.19 6.64 ;
        RECT  103.08 190.585 103.28 191.315 ;
        RECT  103.575 190.585 103.775 191.315 ;
        RECT  104.075 190.585 104.275 191.315 ;
        RECT  104.575 190.585 104.775 191.315 ;
        RECT  105.07 190.585 105.27 191.315 ;
        RECT  105.815 0.17 106.585 0.94 ;
        RECT  105.815 0.17 106.075 12.9 ;
        RECT  106.325 0.17 106.585 12.9 ;
        RECT  105.305 0.52 105.565 5.815 ;
        RECT  105.89 190.585 106.09 191.315 ;
        RECT  106.835 0.17 107.605 0.43 ;
        RECT  106.835 0.17 107.095 11.5 ;
        RECT  107.345 0.17 107.605 11.5 ;
        RECT  106.385 190.585 106.585 191.315 ;
        RECT  106.885 190.585 107.085 191.315 ;
        RECT  107.385 190.585 107.585 191.315 ;
        RECT  108.875 0.17 109.645 0.43 ;
        RECT  108.875 0.17 109.135 10.48 ;
        RECT  109.385 0.17 109.645 10.99 ;
        RECT  107.88 190.585 108.08 191.315 ;
        RECT  108.7 190.585 108.9 191.315 ;
        RECT  109.895 0.17 110.665 0.94 ;
        RECT  109.895 0.17 110.155 8.7 ;
        RECT  110.405 0.17 110.665 12.9 ;
        RECT  109.195 190.585 109.395 191.315 ;
        RECT  109.695 190.585 109.895 191.315 ;
        RECT  110.195 190.585 110.395 191.315 ;
        RECT  110.69 190.585 110.89 191.315 ;
        RECT  110.915 0.52 111.175 2.485 ;
        RECT  111.51 190.585 111.71 191.315 ;
        RECT  111.78 0.52 112.04 14.11 ;
        RECT  112.005 190.585 112.205 191.315 ;
        RECT  112.29 0.52 112.55 2.335 ;
        RECT  112.505 190.585 112.705 191.315 ;
        RECT  113.005 190.585 113.205 191.315 ;
        RECT  113.5 190.585 113.7 191.315 ;
        RECT  115.69 0.52 115.95 5.16 ;
        RECT  115.17 4.9 115.95 5.16 ;
        RECT  115.17 4.9 115.43 6.64 ;
        RECT  114.32 190.585 114.52 191.315 ;
        RECT  114.815 190.585 115.015 191.315 ;
        RECT  115.315 190.585 115.515 191.315 ;
        RECT  115.815 190.585 116.015 191.315 ;
        RECT  116.31 190.585 116.51 191.315 ;
        RECT  117.055 0.17 117.825 0.94 ;
        RECT  117.055 0.17 117.315 12.9 ;
        RECT  117.565 0.17 117.825 12.9 ;
        RECT  116.545 0.52 116.805 5.815 ;
        RECT  117.13 190.585 117.33 191.315 ;
        RECT  118.075 0.17 118.845 0.43 ;
        RECT  118.075 0.17 118.335 11.5 ;
        RECT  118.585 0.17 118.845 11.5 ;
        RECT  117.625 190.585 117.825 191.315 ;
        RECT  118.125 190.585 118.325 191.315 ;
        RECT  118.625 190.585 118.825 191.315 ;
        RECT  120.115 0.17 120.885 0.43 ;
        RECT  120.115 0.17 120.375 10.48 ;
        RECT  120.625 0.17 120.885 10.99 ;
        RECT  119.12 190.585 119.32 191.315 ;
        RECT  119.94 190.585 120.14 191.315 ;
        RECT  121.135 0.17 121.905 0.94 ;
        RECT  121.135 0.17 121.395 8.7 ;
        RECT  121.645 0.17 121.905 12.9 ;
        RECT  120.435 190.585 120.635 191.315 ;
        RECT  120.935 190.585 121.135 191.315 ;
        RECT  121.435 190.585 121.635 191.315 ;
        RECT  121.93 190.585 122.13 191.315 ;
        RECT  122.155 0.52 122.415 2.485 ;
        RECT  122.75 190.585 122.95 191.315 ;
        RECT  123.02 0.52 123.28 14.11 ;
        RECT  123.245 190.585 123.445 191.315 ;
        RECT  123.53 0.52 123.79 2.335 ;
        RECT  123.745 190.585 123.945 191.315 ;
        RECT  124.245 190.585 124.445 191.315 ;
        RECT  124.74 190.585 124.94 191.315 ;
        RECT  126.93 0.52 127.19 5.16 ;
        RECT  126.41 4.9 127.19 5.16 ;
        RECT  126.41 4.9 126.67 6.64 ;
        RECT  125.56 190.585 125.76 191.315 ;
        RECT  126.055 190.585 126.255 191.315 ;
        RECT  126.555 190.585 126.755 191.315 ;
        RECT  127.055 190.585 127.255 191.315 ;
        RECT  127.55 190.585 127.75 191.315 ;
        RECT  128.295 0.17 129.065 0.94 ;
        RECT  128.295 0.17 128.555 12.9 ;
        RECT  128.805 0.17 129.065 12.9 ;
        RECT  127.785 0.52 128.045 5.815 ;
        RECT  128.37 190.585 128.57 191.315 ;
        RECT  129.315 0.17 130.085 0.43 ;
        RECT  129.315 0.17 129.575 11.5 ;
        RECT  129.825 0.17 130.085 11.5 ;
        RECT  128.865 190.585 129.065 191.315 ;
        RECT  129.365 190.585 129.565 191.315 ;
        RECT  129.865 190.585 130.065 191.315 ;
        RECT  131.355 0.17 132.125 0.43 ;
        RECT  131.355 0.17 131.615 10.48 ;
        RECT  131.865 0.17 132.125 10.99 ;
        RECT  130.36 190.585 130.56 191.315 ;
        RECT  131.18 190.585 131.38 191.315 ;
        RECT  132.375 0.17 133.145 0.94 ;
        RECT  132.375 0.17 132.635 8.7 ;
        RECT  132.885 0.17 133.145 12.9 ;
        RECT  131.675 190.585 131.875 191.315 ;
        RECT  132.175 190.585 132.375 191.315 ;
        RECT  132.675 190.585 132.875 191.315 ;
        RECT  133.17 190.585 133.37 191.315 ;
        RECT  133.395 0.52 133.655 2.485 ;
        RECT  133.99 190.585 134.19 191.315 ;
        RECT  134.26 0.52 134.52 14.11 ;
        RECT  134.485 190.585 134.685 191.315 ;
        RECT  134.77 0.52 135.03 2.335 ;
        RECT  134.985 190.585 135.185 191.315 ;
        RECT  135.485 190.585 135.685 191.315 ;
        RECT  135.98 190.585 136.18 191.315 ;
        RECT  138.17 0.52 138.43 5.16 ;
        RECT  137.65 4.9 138.43 5.16 ;
        RECT  137.65 4.9 137.91 6.64 ;
        RECT  136.8 190.585 137 191.315 ;
        RECT  137.295 190.585 137.495 191.315 ;
        RECT  137.795 190.585 137.995 191.315 ;
        RECT  138.295 190.585 138.495 191.315 ;
        RECT  138.79 190.585 138.99 191.315 ;
        RECT  139.535 0.17 140.305 0.94 ;
        RECT  139.535 0.17 139.795 12.9 ;
        RECT  140.045 0.17 140.305 12.9 ;
        RECT  139.025 0.52 139.285 5.815 ;
        RECT  139.61 190.585 139.81 191.315 ;
        RECT  140.555 0.17 141.325 0.43 ;
        RECT  140.555 0.17 140.815 11.5 ;
        RECT  141.065 0.17 141.325 11.5 ;
        RECT  140.105 190.585 140.305 191.315 ;
        RECT  140.605 190.585 140.805 191.315 ;
        RECT  141.105 190.585 141.305 191.315 ;
        RECT  142.595 0.17 143.365 0.43 ;
        RECT  142.595 0.17 142.855 10.48 ;
        RECT  143.105 0.17 143.365 10.99 ;
        RECT  141.6 190.585 141.8 191.315 ;
        RECT  142.42 190.585 142.62 191.315 ;
        RECT  143.615 0.17 144.385 0.94 ;
        RECT  143.615 0.17 143.875 8.7 ;
        RECT  144.125 0.17 144.385 12.9 ;
        RECT  142.915 190.585 143.115 191.315 ;
        RECT  143.415 190.585 143.615 191.315 ;
        RECT  143.915 190.585 144.115 191.315 ;
        RECT  144.41 190.585 144.61 191.315 ;
        RECT  144.635 0.52 144.895 2.485 ;
        RECT  145.23 190.585 145.43 191.315 ;
        RECT  145.5 0.52 145.76 14.11 ;
        RECT  145.725 190.585 145.925 191.315 ;
        RECT  146.01 0.52 146.27 2.335 ;
        RECT  146.225 190.585 146.425 191.315 ;
        RECT  146.725 190.585 146.925 191.315 ;
        RECT  147.22 190.585 147.42 191.315 ;
        RECT  149.41 0.52 149.67 5.16 ;
        RECT  148.89 4.9 149.67 5.16 ;
        RECT  148.89 4.9 149.15 6.64 ;
        RECT  148.04 190.585 148.24 191.315 ;
        RECT  148.535 190.585 148.735 191.315 ;
        RECT  149.035 190.585 149.235 191.315 ;
        RECT  149.535 190.585 149.735 191.315 ;
        RECT  150.03 190.585 150.23 191.315 ;
        RECT  150.775 0.17 151.545 0.94 ;
        RECT  150.775 0.17 151.035 12.9 ;
        RECT  151.285 0.17 151.545 12.9 ;
        RECT  150.265 0.52 150.525 5.815 ;
        RECT  150.85 190.585 151.05 191.315 ;
        RECT  151.795 0.17 152.565 0.43 ;
        RECT  151.795 0.17 152.055 11.5 ;
        RECT  152.305 0.17 152.565 11.5 ;
        RECT  151.345 190.585 151.545 191.315 ;
        RECT  151.845 190.585 152.045 191.315 ;
        RECT  152.345 190.585 152.545 191.315 ;
        RECT  153.835 0.17 154.605 0.43 ;
        RECT  153.835 0.17 154.095 10.48 ;
        RECT  154.345 0.17 154.605 10.99 ;
        RECT  152.84 190.585 153.04 191.315 ;
        RECT  153.66 190.585 153.86 191.315 ;
        RECT  154.855 0.17 155.625 0.94 ;
        RECT  154.855 0.17 155.115 8.7 ;
        RECT  155.365 0.17 155.625 12.9 ;
        RECT  154.155 190.585 154.355 191.315 ;
        RECT  154.655 190.585 154.855 191.315 ;
        RECT  155.155 190.585 155.355 191.315 ;
        RECT  155.65 190.585 155.85 191.315 ;
        RECT  155.875 0.52 156.135 2.485 ;
        RECT  156.47 190.585 156.67 191.315 ;
        RECT  156.74 0.52 157 14.11 ;
        RECT  156.965 190.585 157.165 191.315 ;
        RECT  157.25 0.52 157.51 2.335 ;
        RECT  157.465 190.585 157.665 191.315 ;
        RECT  157.965 190.585 158.165 191.315 ;
        RECT  158.46 190.585 158.66 191.315 ;
        RECT  160.65 0.52 160.91 5.16 ;
        RECT  160.13 4.9 160.91 5.16 ;
        RECT  160.13 4.9 160.39 6.64 ;
        RECT  159.28 190.585 159.48 191.315 ;
        RECT  159.775 190.585 159.975 191.315 ;
        RECT  160.275 190.585 160.475 191.315 ;
        RECT  160.775 190.585 160.975 191.315 ;
        RECT  161.27 190.585 161.47 191.315 ;
        RECT  162.015 0.17 162.785 0.94 ;
        RECT  162.015 0.17 162.275 12.9 ;
        RECT  162.525 0.17 162.785 12.9 ;
        RECT  161.505 0.52 161.765 5.815 ;
        RECT  162.09 190.585 162.29 191.315 ;
        RECT  163.035 0.17 163.805 0.43 ;
        RECT  163.035 0.17 163.295 11.5 ;
        RECT  163.545 0.17 163.805 11.5 ;
        RECT  162.585 190.585 162.785 191.315 ;
        RECT  163.085 190.585 163.285 191.315 ;
        RECT  163.585 190.585 163.785 191.315 ;
        RECT  165.075 0.17 165.845 0.43 ;
        RECT  165.075 0.17 165.335 10.48 ;
        RECT  165.585 0.17 165.845 10.99 ;
        RECT  164.08 190.585 164.28 191.315 ;
        RECT  164.9 190.585 165.1 191.315 ;
        RECT  166.095 0.17 166.865 0.94 ;
        RECT  166.095 0.17 166.355 8.7 ;
        RECT  166.605 0.17 166.865 12.9 ;
        RECT  165.395 190.585 165.595 191.315 ;
        RECT  165.895 190.585 166.095 191.315 ;
        RECT  166.395 190.585 166.595 191.315 ;
        RECT  166.89 190.585 167.09 191.315 ;
        RECT  167.115 0.52 167.375 2.485 ;
        RECT  167.71 190.585 167.91 191.315 ;
        RECT  167.98 0.52 168.24 14.11 ;
        RECT  168.205 190.585 168.405 191.315 ;
        RECT  168.49 0.52 168.75 2.335 ;
        RECT  168.705 190.585 168.905 191.315 ;
        RECT  169.205 190.585 169.405 191.315 ;
        RECT  169.7 190.585 169.9 191.315 ;
        RECT  171.89 0.52 172.15 5.16 ;
        RECT  171.37 4.9 172.15 5.16 ;
        RECT  171.37 4.9 171.63 6.64 ;
        RECT  170.52 190.585 170.72 191.315 ;
        RECT  171.015 190.585 171.215 191.315 ;
        RECT  171.515 190.585 171.715 191.315 ;
        RECT  172.015 190.585 172.215 191.315 ;
        RECT  172.51 190.585 172.71 191.315 ;
        RECT  173.255 0.17 174.025 0.94 ;
        RECT  173.255 0.17 173.515 12.9 ;
        RECT  173.765 0.17 174.025 12.9 ;
        RECT  172.745 0.52 173.005 5.815 ;
        RECT  173.33 190.585 173.53 191.315 ;
        RECT  174.275 0.17 175.045 0.43 ;
        RECT  174.275 0.17 174.535 11.5 ;
        RECT  174.785 0.17 175.045 11.5 ;
        RECT  173.825 190.585 174.025 191.315 ;
        RECT  174.325 190.585 174.525 191.315 ;
        RECT  174.825 190.585 175.025 191.315 ;
        RECT  176.315 0.17 177.085 0.43 ;
        RECT  176.315 0.17 176.575 10.48 ;
        RECT  176.825 0.17 177.085 10.99 ;
        RECT  175.32 190.585 175.52 191.315 ;
        RECT  176.14 190.585 176.34 191.315 ;
        RECT  177.335 0.17 178.105 0.94 ;
        RECT  177.335 0.17 177.595 8.7 ;
        RECT  177.845 0.17 178.105 12.9 ;
        RECT  176.635 190.585 176.835 191.315 ;
        RECT  177.135 190.585 177.335 191.315 ;
        RECT  177.635 190.585 177.835 191.315 ;
        RECT  178.13 190.585 178.33 191.315 ;
        RECT  178.355 0.52 178.615 2.485 ;
        RECT  178.95 190.585 179.15 191.315 ;
        RECT  179.22 0.52 179.48 14.11 ;
        RECT  179.445 190.585 179.645 191.315 ;
        RECT  179.73 0.52 179.99 2.335 ;
        RECT  179.945 190.585 180.145 191.315 ;
        RECT  180.445 190.585 180.645 191.315 ;
        RECT  180.94 190.585 181.14 191.315 ;
        RECT  183.13 0.52 183.39 5.16 ;
        RECT  182.61 4.9 183.39 5.16 ;
        RECT  182.61 4.9 182.87 6.64 ;
        RECT  181.76 190.585 181.96 191.315 ;
        RECT  182.255 190.585 182.455 191.315 ;
        RECT  182.755 190.585 182.955 191.315 ;
        RECT  183.255 190.585 183.455 191.315 ;
        RECT  183.75 190.585 183.95 191.315 ;
        RECT  184.495 0.17 185.265 0.94 ;
        RECT  184.495 0.17 184.755 12.9 ;
        RECT  185.005 0.17 185.265 12.9 ;
        RECT  183.985 0.52 184.245 5.815 ;
        RECT  184.57 190.585 184.77 191.315 ;
        RECT  185.515 0.17 186.285 0.43 ;
        RECT  185.515 0.17 185.775 11.5 ;
        RECT  186.025 0.17 186.285 11.5 ;
        RECT  185.065 190.585 185.265 191.315 ;
        RECT  185.565 190.585 185.765 191.315 ;
        RECT  186.065 190.585 186.265 191.315 ;
        RECT  187.555 0.17 188.325 0.43 ;
        RECT  187.555 0.17 187.815 10.48 ;
        RECT  188.065 0.17 188.325 10.99 ;
        RECT  186.56 190.585 186.76 191.315 ;
        RECT  187.38 190.585 187.58 191.315 ;
        RECT  188.575 0.17 189.345 0.94 ;
        RECT  188.575 0.17 188.835 8.7 ;
        RECT  189.085 0.17 189.345 12.9 ;
        RECT  187.875 190.585 188.075 191.315 ;
        RECT  188.375 190.585 188.575 191.315 ;
        RECT  188.875 190.585 189.075 191.315 ;
        RECT  189.37 190.585 189.57 191.315 ;
        RECT  189.595 0.52 189.855 2.485 ;
        RECT  190.19 190.585 190.39 191.315 ;
        RECT  190.46 0.52 190.72 14.11 ;
        RECT  190.685 190.585 190.885 191.315 ;
        RECT  190.97 0.52 191.23 2.335 ;
        RECT  191.185 190.585 191.385 191.315 ;
        RECT  191.685 190.585 191.885 191.315 ;
        RECT  192.18 190.585 192.38 191.315 ;
        RECT  194.37 0.52 194.63 5.16 ;
        RECT  193.85 4.9 194.63 5.16 ;
        RECT  193.85 4.9 194.11 6.64 ;
        RECT  193 190.585 193.2 191.315 ;
        RECT  193.495 190.585 193.695 191.315 ;
        RECT  193.995 190.585 194.195 191.315 ;
        RECT  194.495 190.585 194.695 191.315 ;
        RECT  194.99 190.585 195.19 191.315 ;
        RECT  195.735 0.17 196.505 0.94 ;
        RECT  195.735 0.17 195.995 12.9 ;
        RECT  196.245 0.17 196.505 12.9 ;
        RECT  195.225 0.52 195.485 5.815 ;
        RECT  195.81 190.585 196.01 191.315 ;
        RECT  196.755 0.17 197.525 0.43 ;
        RECT  196.755 0.17 197.015 11.5 ;
        RECT  197.265 0.17 197.525 11.5 ;
        RECT  196.305 190.585 196.505 191.315 ;
        RECT  196.805 190.585 197.005 191.315 ;
        RECT  197.305 190.585 197.505 191.315 ;
        RECT  198.795 0.17 199.565 0.43 ;
        RECT  198.795 0.17 199.055 10.48 ;
        RECT  199.305 0.17 199.565 10.99 ;
        RECT  197.8 190.585 198 191.315 ;
        RECT  198.62 190.585 198.82 191.315 ;
        RECT  199.815 0.17 200.585 0.94 ;
        RECT  199.815 0.17 200.075 8.7 ;
        RECT  200.325 0.17 200.585 12.9 ;
        RECT  199.115 190.585 199.315 191.315 ;
        RECT  199.615 190.585 199.815 191.315 ;
        RECT  200.115 190.585 200.315 191.315 ;
        RECT  200.61 190.585 200.81 191.315 ;
        RECT  200.835 0.52 201.095 2.485 ;
        RECT  201.43 190.585 201.63 191.315 ;
        RECT  201.7 0.52 201.96 14.11 ;
        RECT  201.925 190.585 202.125 191.315 ;
        RECT  202.21 0.52 202.47 2.335 ;
        RECT  202.425 190.585 202.625 191.315 ;
        RECT  202.925 190.585 203.125 191.315 ;
        RECT  203.42 190.585 203.62 191.315 ;
        RECT  205.61 0.52 205.87 5.16 ;
        RECT  205.09 4.9 205.87 5.16 ;
        RECT  205.09 4.9 205.35 6.64 ;
        RECT  204.24 190.585 204.44 191.315 ;
        RECT  204.735 190.585 204.935 191.315 ;
        RECT  205.235 190.585 205.435 191.315 ;
        RECT  205.735 190.585 205.935 191.315 ;
        RECT  206.23 190.585 206.43 191.315 ;
        RECT  206.975 0.17 207.745 0.94 ;
        RECT  206.975 0.17 207.235 12.9 ;
        RECT  207.485 0.17 207.745 12.9 ;
        RECT  206.465 0.52 206.725 5.815 ;
        RECT  207.05 190.585 207.25 191.315 ;
        RECT  207.995 0.17 208.765 0.43 ;
        RECT  207.995 0.17 208.255 11.5 ;
        RECT  208.505 0.17 208.765 11.5 ;
        RECT  207.545 190.585 207.745 191.315 ;
        RECT  208.045 190.585 208.245 191.315 ;
        RECT  208.545 190.585 208.745 191.315 ;
        RECT  210.035 0.17 210.805 0.43 ;
        RECT  210.035 0.17 210.295 10.48 ;
        RECT  210.545 0.17 210.805 10.99 ;
        RECT  209.04 190.585 209.24 191.315 ;
        RECT  209.86 190.585 210.06 191.315 ;
        RECT  211.055 0.17 211.825 0.94 ;
        RECT  211.055 0.17 211.315 8.7 ;
        RECT  211.565 0.17 211.825 12.9 ;
        RECT  210.355 190.585 210.555 191.315 ;
        RECT  210.855 190.585 211.055 191.315 ;
        RECT  211.355 190.585 211.555 191.315 ;
        RECT  211.85 190.585 212.05 191.315 ;
        RECT  212.075 0.52 212.335 2.485 ;
        RECT  212.67 190.585 212.87 191.315 ;
        RECT  212.94 0.52 213.2 14.11 ;
        RECT  213.165 190.585 213.365 191.315 ;
        RECT  213.45 0.52 213.71 2.335 ;
        RECT  213.665 190.585 213.865 191.315 ;
        RECT  214.165 190.585 214.365 191.315 ;
        RECT  214.66 190.585 214.86 191.315 ;
        RECT  216.85 0.52 217.11 5.16 ;
        RECT  216.33 4.9 217.11 5.16 ;
        RECT  216.33 4.9 216.59 6.64 ;
        RECT  215.48 190.585 215.68 191.315 ;
        RECT  215.975 190.585 216.175 191.315 ;
        RECT  216.475 190.585 216.675 191.315 ;
        RECT  216.975 190.585 217.175 191.315 ;
        RECT  217.47 190.585 217.67 191.315 ;
        RECT  218.215 0.17 218.985 0.94 ;
        RECT  218.215 0.17 218.475 12.9 ;
        RECT  218.725 0.17 218.985 12.9 ;
        RECT  217.705 0.52 217.965 5.815 ;
        RECT  218.29 190.585 218.49 191.315 ;
        RECT  219.235 0.17 220.005 0.43 ;
        RECT  219.235 0.17 219.495 11.5 ;
        RECT  219.745 0.17 220.005 11.5 ;
        RECT  218.785 190.585 218.985 191.315 ;
        RECT  219.285 190.585 219.485 191.315 ;
        RECT  219.785 190.585 219.985 191.315 ;
        RECT  221.275 0.17 222.045 0.43 ;
        RECT  221.275 0.17 221.535 10.48 ;
        RECT  221.785 0.17 222.045 10.99 ;
        RECT  220.28 190.585 220.48 191.315 ;
        RECT  221.1 190.585 221.3 191.315 ;
        RECT  222.295 0.17 223.065 0.94 ;
        RECT  222.295 0.17 222.555 8.7 ;
        RECT  222.805 0.17 223.065 12.9 ;
        RECT  221.595 190.585 221.795 191.315 ;
        RECT  222.095 190.585 222.295 191.315 ;
        RECT  222.595 190.585 222.795 191.315 ;
        RECT  223.09 190.585 223.29 191.315 ;
        RECT  223.315 0.52 223.575 2.485 ;
        RECT  223.91 190.585 224.11 191.315 ;
        RECT  224.18 0.52 224.44 14.11 ;
        RECT  224.405 190.585 224.605 191.315 ;
        RECT  224.69 0.52 224.95 2.335 ;
        RECT  224.905 190.585 225.105 191.315 ;
        RECT  225.405 190.585 225.605 191.315 ;
        RECT  225.9 190.585 226.1 191.315 ;
        RECT  228.09 0.52 228.35 5.16 ;
        RECT  227.57 4.9 228.35 5.16 ;
        RECT  227.57 4.9 227.83 6.64 ;
        RECT  226.72 190.585 226.92 191.315 ;
        RECT  227.215 190.585 227.415 191.315 ;
        RECT  227.715 190.585 227.915 191.315 ;
        RECT  228.215 190.585 228.415 191.315 ;
        RECT  228.71 190.585 228.91 191.315 ;
        RECT  229.455 0.17 230.225 0.94 ;
        RECT  229.455 0.17 229.715 12.9 ;
        RECT  229.965 0.17 230.225 12.9 ;
        RECT  228.945 0.52 229.205 5.815 ;
        RECT  229.53 190.585 229.73 191.315 ;
        RECT  230.475 0.17 231.245 0.43 ;
        RECT  230.475 0.17 230.735 11.5 ;
        RECT  230.985 0.17 231.245 11.5 ;
        RECT  230.025 190.585 230.225 191.315 ;
        RECT  230.525 190.585 230.725 191.315 ;
        RECT  231.025 190.585 231.225 191.315 ;
        RECT  232.515 0.17 233.285 0.43 ;
        RECT  232.515 0.17 232.775 10.48 ;
        RECT  233.025 0.17 233.285 10.99 ;
        RECT  231.52 190.585 231.72 191.315 ;
        RECT  232.34 190.585 232.54 191.315 ;
        RECT  233.535 0.17 234.305 0.94 ;
        RECT  233.535 0.17 233.795 8.7 ;
        RECT  234.045 0.17 234.305 12.9 ;
        RECT  232.835 190.585 233.035 191.315 ;
        RECT  233.335 190.585 233.535 191.315 ;
        RECT  233.835 190.585 234.035 191.315 ;
        RECT  234.33 190.585 234.53 191.315 ;
        RECT  234.555 0.52 234.815 2.485 ;
        RECT  235.15 190.585 235.35 191.315 ;
        RECT  235.42 0.52 235.68 14.11 ;
        RECT  235.645 190.585 235.845 191.315 ;
        RECT  235.93 0.52 236.19 2.335 ;
        RECT  236.145 190.585 236.345 191.315 ;
        RECT  236.645 190.585 236.845 191.315 ;
        RECT  237.14 190.585 237.34 191.315 ;
        RECT  239.33 0.52 239.59 5.16 ;
        RECT  238.81 4.9 239.59 5.16 ;
        RECT  238.81 4.9 239.07 6.64 ;
        RECT  237.96 190.585 238.16 191.315 ;
        RECT  238.455 190.585 238.655 191.315 ;
        RECT  238.955 190.585 239.155 191.315 ;
        RECT  239.455 190.585 239.655 191.315 ;
        RECT  239.95 190.585 240.15 191.315 ;
        RECT  240.695 0.17 241.465 0.94 ;
        RECT  240.695 0.17 240.955 12.9 ;
        RECT  241.205 0.17 241.465 12.9 ;
        RECT  240.185 0.52 240.445 5.815 ;
        RECT  240.77 190.585 240.97 191.315 ;
        RECT  241.715 0.17 242.485 0.43 ;
        RECT  241.715 0.17 241.975 11.5 ;
        RECT  242.225 0.17 242.485 11.5 ;
        RECT  241.265 190.585 241.465 191.315 ;
        RECT  241.765 190.585 241.965 191.315 ;
        RECT  242.265 190.585 242.465 191.315 ;
        RECT  243.755 0.17 244.525 0.43 ;
        RECT  243.755 0.17 244.015 10.48 ;
        RECT  244.265 0.17 244.525 10.99 ;
        RECT  242.76 190.585 242.96 191.315 ;
        RECT  243.58 190.585 243.78 191.315 ;
        RECT  244.775 0.17 245.545 0.94 ;
        RECT  244.775 0.17 245.035 8.7 ;
        RECT  245.285 0.17 245.545 12.9 ;
        RECT  244.075 190.585 244.275 191.315 ;
        RECT  244.575 190.585 244.775 191.315 ;
        RECT  245.075 190.585 245.275 191.315 ;
        RECT  245.57 190.585 245.77 191.315 ;
        RECT  245.795 0.52 246.055 2.485 ;
        RECT  246.39 190.585 246.59 191.315 ;
        RECT  246.66 0.52 246.92 14.11 ;
        RECT  246.885 190.585 247.085 191.315 ;
        RECT  247.17 0.52 247.43 2.335 ;
        RECT  247.385 190.585 247.585 191.315 ;
        RECT  247.885 190.585 248.085 191.315 ;
        RECT  248.38 190.585 248.58 191.315 ;
        RECT  250.57 0.52 250.83 5.16 ;
        RECT  250.05 4.9 250.83 5.16 ;
        RECT  250.05 4.9 250.31 6.64 ;
        RECT  249.2 190.585 249.4 191.315 ;
        RECT  249.695 190.585 249.895 191.315 ;
        RECT  250.195 190.585 250.395 191.315 ;
        RECT  250.695 190.585 250.895 191.315 ;
        RECT  251.19 190.585 251.39 191.315 ;
        RECT  251.935 0.17 252.705 0.94 ;
        RECT  251.935 0.17 252.195 12.9 ;
        RECT  252.445 0.17 252.705 12.9 ;
        RECT  251.425 0.52 251.685 5.815 ;
        RECT  252.01 190.585 252.21 191.315 ;
        RECT  252.955 0.17 253.725 0.43 ;
        RECT  252.955 0.17 253.215 11.5 ;
        RECT  253.465 0.17 253.725 11.5 ;
        RECT  252.505 190.585 252.705 191.315 ;
        RECT  253.005 190.585 253.205 191.315 ;
        RECT  253.505 190.585 253.705 191.315 ;
        RECT  254.995 0.17 255.765 0.43 ;
        RECT  254.995 0.17 255.255 10.48 ;
        RECT  255.505 0.17 255.765 10.99 ;
        RECT  254 190.585 254.2 191.315 ;
        RECT  254.82 190.585 255.02 191.315 ;
        RECT  256.015 0.17 256.785 0.94 ;
        RECT  256.015 0.17 256.275 8.7 ;
        RECT  256.525 0.17 256.785 12.9 ;
        RECT  255.315 190.585 255.515 191.315 ;
        RECT  255.815 190.585 256.015 191.315 ;
        RECT  256.315 190.585 256.515 191.315 ;
        RECT  256.81 190.585 257.01 191.315 ;
        RECT  257.035 0.52 257.295 2.485 ;
        RECT  257.63 190.585 257.83 191.315 ;
        RECT  257.9 0.52 258.16 14.11 ;
        RECT  258.125 190.585 258.325 191.315 ;
        RECT  258.41 0.52 258.67 2.335 ;
        RECT  258.625 190.585 258.825 191.315 ;
        RECT  259.125 190.585 259.325 191.315 ;
        RECT  259.62 190.585 259.82 191.315 ;
        RECT  261.81 0.52 262.07 5.16 ;
        RECT  261.29 4.9 262.07 5.16 ;
        RECT  261.29 4.9 261.55 6.64 ;
        RECT  260.44 190.585 260.64 191.315 ;
        RECT  260.935 190.585 261.135 191.315 ;
        RECT  261.435 190.585 261.635 191.315 ;
        RECT  261.935 190.585 262.135 191.315 ;
        RECT  262.43 190.585 262.63 191.315 ;
        RECT  263.175 0.17 263.945 0.94 ;
        RECT  263.175 0.17 263.435 12.9 ;
        RECT  263.685 0.17 263.945 12.9 ;
        RECT  262.665 0.52 262.925 5.815 ;
        RECT  263.25 190.585 263.45 191.315 ;
        RECT  264.195 0.17 264.965 0.43 ;
        RECT  264.195 0.17 264.455 11.5 ;
        RECT  264.705 0.17 264.965 11.5 ;
        RECT  263.745 190.585 263.945 191.315 ;
        RECT  264.245 190.585 264.445 191.315 ;
        RECT  264.745 190.585 264.945 191.315 ;
        RECT  266.235 0.17 267.005 0.43 ;
        RECT  266.235 0.17 266.495 10.48 ;
        RECT  266.745 0.17 267.005 10.99 ;
        RECT  265.24 190.585 265.44 191.315 ;
        RECT  266.06 190.585 266.26 191.315 ;
        RECT  267.255 0.17 268.025 0.94 ;
        RECT  267.255 0.17 267.515 8.7 ;
        RECT  267.765 0.17 268.025 12.9 ;
        RECT  266.555 190.585 266.755 191.315 ;
        RECT  267.055 190.585 267.255 191.315 ;
        RECT  267.555 190.585 267.755 191.315 ;
        RECT  268.05 190.585 268.25 191.315 ;
        RECT  268.275 0.52 268.535 2.485 ;
        RECT  268.87 190.585 269.07 191.315 ;
        RECT  269.14 0.52 269.4 14.11 ;
        RECT  269.365 190.585 269.565 191.315 ;
        RECT  269.65 0.52 269.91 2.335 ;
        RECT  269.865 190.585 270.065 191.315 ;
        RECT  270.365 190.585 270.565 191.315 ;
        RECT  270.86 190.585 271.06 191.315 ;
        RECT  273.05 0.52 273.31 5.16 ;
        RECT  272.53 4.9 273.31 5.16 ;
        RECT  272.53 4.9 272.79 6.64 ;
        RECT  271.68 190.585 271.88 191.315 ;
        RECT  272.175 190.585 272.375 191.315 ;
        RECT  272.675 190.585 272.875 191.315 ;
        RECT  273.175 190.585 273.375 191.315 ;
        RECT  273.67 190.585 273.87 191.315 ;
        RECT  274.415 0.17 275.185 0.94 ;
        RECT  274.415 0.17 274.675 12.9 ;
        RECT  274.925 0.17 275.185 12.9 ;
        RECT  273.905 0.52 274.165 5.815 ;
        RECT  274.49 190.585 274.69 191.315 ;
        RECT  275.435 0.17 276.205 0.43 ;
        RECT  275.435 0.17 275.695 11.5 ;
        RECT  275.945 0.17 276.205 11.5 ;
        RECT  274.985 190.585 275.185 191.315 ;
        RECT  275.485 190.585 275.685 191.315 ;
        RECT  275.985 190.585 276.185 191.315 ;
        RECT  277.475 0.17 278.245 0.43 ;
        RECT  277.475 0.17 277.735 10.48 ;
        RECT  277.985 0.17 278.245 10.99 ;
        RECT  276.48 190.585 276.68 191.315 ;
        RECT  277.3 190.585 277.5 191.315 ;
        RECT  278.495 0.17 279.265 0.94 ;
        RECT  278.495 0.17 278.755 8.7 ;
        RECT  279.005 0.17 279.265 12.9 ;
        RECT  277.795 190.585 277.995 191.315 ;
        RECT  278.295 190.585 278.495 191.315 ;
        RECT  278.795 190.585 278.995 191.315 ;
        RECT  279.29 190.585 279.49 191.315 ;
        RECT  279.515 0.52 279.775 2.485 ;
        RECT  280.11 190.585 280.31 191.315 ;
        RECT  280.38 0.52 280.64 14.11 ;
        RECT  280.605 190.585 280.805 191.315 ;
        RECT  280.89 0.52 281.15 2.335 ;
        RECT  281.105 190.585 281.305 191.315 ;
        RECT  281.605 190.585 281.805 191.315 ;
        RECT  282.1 190.585 282.3 191.315 ;
        RECT  284.29 0.52 284.55 5.16 ;
        RECT  283.77 4.9 284.55 5.16 ;
        RECT  283.77 4.9 284.03 6.64 ;
        RECT  282.92 190.585 283.12 191.315 ;
        RECT  283.415 190.585 283.615 191.315 ;
        RECT  283.915 190.585 284.115 191.315 ;
        RECT  284.415 190.585 284.615 191.315 ;
        RECT  284.91 190.585 285.11 191.315 ;
        RECT  285.655 0.17 286.425 0.94 ;
        RECT  285.655 0.17 285.915 12.9 ;
        RECT  286.165 0.17 286.425 12.9 ;
        RECT  285.145 0.52 285.405 5.815 ;
        RECT  285.73 190.585 285.93 191.315 ;
        RECT  286.675 0.17 287.445 0.43 ;
        RECT  286.675 0.17 286.935 11.5 ;
        RECT  287.185 0.17 287.445 11.5 ;
        RECT  286.225 190.585 286.425 191.315 ;
        RECT  286.725 190.585 286.925 191.315 ;
        RECT  287.225 190.585 287.425 191.315 ;
        RECT  288.715 0.17 289.485 0.43 ;
        RECT  288.715 0.17 288.975 10.48 ;
        RECT  289.225 0.17 289.485 10.99 ;
        RECT  287.72 190.585 287.92 191.315 ;
        RECT  288.54 190.585 288.74 191.315 ;
        RECT  289.735 0.17 290.505 0.94 ;
        RECT  289.735 0.17 289.995 8.7 ;
        RECT  290.245 0.17 290.505 12.9 ;
        RECT  289.035 190.585 289.235 191.315 ;
        RECT  289.535 190.585 289.735 191.315 ;
        RECT  290.035 190.585 290.235 191.315 ;
        RECT  290.53 190.585 290.73 191.315 ;
        RECT  290.755 0.52 291.015 2.485 ;
        RECT  291.35 190.585 291.55 191.315 ;
        RECT  291.62 0.52 291.88 14.11 ;
        RECT  291.845 190.585 292.045 191.315 ;
        RECT  292.13 0.52 292.39 2.335 ;
        RECT  292.345 190.585 292.545 191.315 ;
        RECT  292.845 190.585 293.045 191.315 ;
        RECT  293.34 190.585 293.54 191.315 ;
        RECT  295.53 0.52 295.79 5.16 ;
        RECT  295.01 4.9 295.79 5.16 ;
        RECT  295.01 4.9 295.27 6.64 ;
        RECT  294.16 190.585 294.36 191.315 ;
        RECT  294.655 190.585 294.855 191.315 ;
        RECT  295.155 190.585 295.355 191.315 ;
        RECT  295.655 190.585 295.855 191.315 ;
        RECT  296.15 190.585 296.35 191.315 ;
        RECT  296.895 0.17 297.665 0.94 ;
        RECT  296.895 0.17 297.155 12.9 ;
        RECT  297.405 0.17 297.665 12.9 ;
        RECT  296.385 0.52 296.645 5.815 ;
        RECT  296.97 190.585 297.17 191.315 ;
        RECT  297.915 0.17 298.685 0.43 ;
        RECT  297.915 0.17 298.175 11.5 ;
        RECT  298.425 0.17 298.685 11.5 ;
        RECT  297.465 190.585 297.665 191.315 ;
        RECT  297.965 190.585 298.165 191.315 ;
        RECT  298.465 190.585 298.665 191.315 ;
        RECT  299.955 0.17 300.725 0.43 ;
        RECT  299.955 0.17 300.215 10.48 ;
        RECT  300.465 0.17 300.725 10.99 ;
        RECT  298.96 190.585 299.16 191.315 ;
        RECT  299.78 190.585 299.98 191.315 ;
        RECT  300.975 0.17 301.745 0.94 ;
        RECT  300.975 0.17 301.235 8.7 ;
        RECT  301.485 0.17 301.745 12.9 ;
        RECT  300.275 190.585 300.475 191.315 ;
        RECT  300.775 190.585 300.975 191.315 ;
        RECT  301.275 190.585 301.475 191.315 ;
        RECT  301.77 190.585 301.97 191.315 ;
        RECT  301.995 0.52 302.255 2.485 ;
        RECT  302.59 190.585 302.79 191.315 ;
        RECT  302.86 0.52 303.12 14.11 ;
        RECT  303.085 190.585 303.285 191.315 ;
        RECT  303.37 0.52 303.63 2.335 ;
        RECT  303.585 190.585 303.785 191.315 ;
        RECT  304.085 190.585 304.285 191.315 ;
        RECT  304.58 190.585 304.78 191.315 ;
        RECT  306.77 0.52 307.03 5.16 ;
        RECT  306.25 4.9 307.03 5.16 ;
        RECT  306.25 4.9 306.51 6.64 ;
        RECT  305.4 190.585 305.6 191.315 ;
        RECT  305.895 190.585 306.095 191.315 ;
        RECT  306.395 190.585 306.595 191.315 ;
        RECT  306.895 190.585 307.095 191.315 ;
        RECT  307.39 190.585 307.59 191.315 ;
        RECT  308.135 0.17 308.905 0.94 ;
        RECT  308.135 0.17 308.395 12.9 ;
        RECT  308.645 0.17 308.905 12.9 ;
        RECT  307.625 0.52 307.885 5.815 ;
        RECT  308.21 190.585 308.41 191.315 ;
        RECT  309.155 0.17 309.925 0.43 ;
        RECT  309.155 0.17 309.415 11.5 ;
        RECT  309.665 0.17 309.925 11.5 ;
        RECT  308.705 190.585 308.905 191.315 ;
        RECT  309.205 190.585 309.405 191.315 ;
        RECT  309.705 190.585 309.905 191.315 ;
        RECT  311.195 0.17 311.965 0.43 ;
        RECT  311.195 0.17 311.455 10.48 ;
        RECT  311.705 0.17 311.965 10.99 ;
        RECT  310.2 190.585 310.4 191.315 ;
        RECT  311.02 190.585 311.22 191.315 ;
        RECT  312.215 0.17 312.985 0.94 ;
        RECT  312.215 0.17 312.475 8.7 ;
        RECT  312.725 0.17 312.985 12.9 ;
        RECT  311.515 190.585 311.715 191.315 ;
        RECT  312.015 190.585 312.215 191.315 ;
        RECT  312.515 190.585 312.715 191.315 ;
        RECT  313.01 190.585 313.21 191.315 ;
        RECT  313.235 0.52 313.495 2.485 ;
        RECT  313.83 190.585 314.03 191.315 ;
        RECT  314.1 0.52 314.36 14.11 ;
        RECT  314.325 190.585 314.525 191.315 ;
        RECT  314.61 0.52 314.87 2.335 ;
        RECT  314.825 190.585 315.025 191.315 ;
        RECT  315.325 190.585 315.525 191.315 ;
        RECT  315.82 190.585 316.02 191.315 ;
        RECT  318.01 0.52 318.27 5.16 ;
        RECT  317.49 4.9 318.27 5.16 ;
        RECT  317.49 4.9 317.75 6.64 ;
        RECT  316.64 190.585 316.84 191.315 ;
        RECT  317.135 190.585 317.335 191.315 ;
        RECT  317.635 190.585 317.835 191.315 ;
        RECT  318.135 190.585 318.335 191.315 ;
        RECT  318.63 190.585 318.83 191.315 ;
        RECT  319.375 0.17 320.145 0.94 ;
        RECT  319.375 0.17 319.635 12.9 ;
        RECT  319.885 0.17 320.145 12.9 ;
        RECT  318.865 0.52 319.125 5.815 ;
        RECT  319.45 190.585 319.65 191.315 ;
        RECT  320.395 0.17 321.165 0.43 ;
        RECT  320.395 0.17 320.655 11.5 ;
        RECT  320.905 0.17 321.165 11.5 ;
        RECT  319.945 190.585 320.145 191.315 ;
        RECT  320.445 190.585 320.645 191.315 ;
        RECT  320.945 190.585 321.145 191.315 ;
        RECT  322.435 0.17 323.205 0.43 ;
        RECT  322.435 0.17 322.695 10.48 ;
        RECT  322.945 0.17 323.205 10.99 ;
        RECT  321.44 190.585 321.64 191.315 ;
        RECT  322.26 190.585 322.46 191.315 ;
        RECT  323.455 0.17 324.225 0.94 ;
        RECT  323.455 0.17 323.715 8.7 ;
        RECT  323.965 0.17 324.225 12.9 ;
        RECT  322.755 190.585 322.955 191.315 ;
        RECT  323.255 190.585 323.455 191.315 ;
        RECT  323.755 190.585 323.955 191.315 ;
        RECT  324.25 190.585 324.45 191.315 ;
        RECT  324.475 0.52 324.735 2.485 ;
        RECT  325.07 190.585 325.27 191.315 ;
        RECT  325.34 0.52 325.6 14.11 ;
        RECT  325.565 190.585 325.765 191.315 ;
        RECT  325.85 0.52 326.11 2.335 ;
        RECT  326.065 190.585 326.265 191.315 ;
        RECT  326.565 190.585 326.765 191.315 ;
        RECT  327.06 190.585 327.26 191.315 ;
        RECT  329.25 0.52 329.51 5.16 ;
        RECT  328.73 4.9 329.51 5.16 ;
        RECT  328.73 4.9 328.99 6.64 ;
        RECT  327.88 190.585 328.08 191.315 ;
        RECT  328.375 190.585 328.575 191.315 ;
        RECT  328.875 190.585 329.075 191.315 ;
        RECT  329.375 190.585 329.575 191.315 ;
        RECT  329.87 190.585 330.07 191.315 ;
        RECT  330.615 0.17 331.385 0.94 ;
        RECT  330.615 0.17 330.875 12.9 ;
        RECT  331.125 0.17 331.385 12.9 ;
        RECT  330.105 0.52 330.365 5.815 ;
        RECT  330.69 190.585 330.89 191.315 ;
        RECT  331.635 0.17 332.405 0.43 ;
        RECT  331.635 0.17 331.895 11.5 ;
        RECT  332.145 0.17 332.405 11.5 ;
        RECT  331.185 190.585 331.385 191.315 ;
        RECT  331.685 190.585 331.885 191.315 ;
        RECT  332.185 190.585 332.385 191.315 ;
        RECT  333.675 0.17 334.445 0.43 ;
        RECT  333.675 0.17 333.935 10.48 ;
        RECT  334.185 0.17 334.445 10.99 ;
        RECT  332.68 190.585 332.88 191.315 ;
        RECT  333.5 190.585 333.7 191.315 ;
        RECT  334.695 0.17 335.465 0.94 ;
        RECT  334.695 0.17 334.955 8.7 ;
        RECT  335.205 0.17 335.465 12.9 ;
        RECT  333.995 190.585 334.195 191.315 ;
        RECT  334.495 190.585 334.695 191.315 ;
        RECT  334.995 190.585 335.195 191.315 ;
        RECT  335.49 190.585 335.69 191.315 ;
        RECT  335.715 0.52 335.975 2.485 ;
        RECT  336.31 190.585 336.51 191.315 ;
        RECT  336.58 0.52 336.84 14.11 ;
        RECT  336.805 190.585 337.005 191.315 ;
        RECT  337.09 0.52 337.35 2.335 ;
        RECT  337.305 190.585 337.505 191.315 ;
        RECT  337.805 190.585 338.005 191.315 ;
        RECT  338.3 190.585 338.5 191.315 ;
        RECT  340.49 0.52 340.75 5.16 ;
        RECT  339.97 4.9 340.75 5.16 ;
        RECT  339.97 4.9 340.23 6.64 ;
        RECT  339.12 190.585 339.32 191.315 ;
        RECT  339.615 190.585 339.815 191.315 ;
        RECT  340.115 190.585 340.315 191.315 ;
        RECT  340.615 190.585 340.815 191.315 ;
        RECT  341.11 190.585 341.31 191.315 ;
        RECT  341.855 0.17 342.625 0.94 ;
        RECT  341.855 0.17 342.115 12.9 ;
        RECT  342.365 0.17 342.625 12.9 ;
        RECT  341.345 0.52 341.605 5.815 ;
        RECT  341.93 190.585 342.13 191.315 ;
        RECT  342.875 0.17 343.645 0.43 ;
        RECT  342.875 0.17 343.135 11.5 ;
        RECT  343.385 0.17 343.645 11.5 ;
        RECT  342.425 190.585 342.625 191.315 ;
        RECT  342.925 190.585 343.125 191.315 ;
        RECT  343.425 190.585 343.625 191.315 ;
        RECT  344.915 0.17 345.685 0.43 ;
        RECT  344.915 0.17 345.175 10.48 ;
        RECT  345.425 0.17 345.685 10.99 ;
        RECT  343.92 190.585 344.12 191.315 ;
        RECT  344.74 190.585 344.94 191.315 ;
        RECT  345.935 0.17 346.705 0.94 ;
        RECT  345.935 0.17 346.195 8.7 ;
        RECT  346.445 0.17 346.705 12.9 ;
        RECT  345.235 190.585 345.435 191.315 ;
        RECT  345.735 190.585 345.935 191.315 ;
        RECT  346.235 190.585 346.435 191.315 ;
        RECT  346.73 190.585 346.93 191.315 ;
        RECT  346.955 0.52 347.215 2.485 ;
        RECT  347.55 190.585 347.75 191.315 ;
        RECT  347.82 0.52 348.08 14.11 ;
        RECT  348.045 190.585 348.245 191.315 ;
        RECT  348.33 0.52 348.59 2.335 ;
        RECT  348.545 190.585 348.745 191.315 ;
        RECT  349.045 190.585 349.245 191.315 ;
        RECT  349.54 190.585 349.74 191.315 ;
        RECT  351.73 0.52 351.99 5.16 ;
        RECT  351.21 4.9 351.99 5.16 ;
        RECT  351.21 4.9 351.47 6.64 ;
        RECT  350.36 190.585 350.56 191.315 ;
        RECT  350.855 190.585 351.055 191.315 ;
        RECT  351.355 190.585 351.555 191.315 ;
        RECT  351.855 190.585 352.055 191.315 ;
        RECT  352.35 190.585 352.55 191.315 ;
        RECT  353.095 0.17 353.865 0.94 ;
        RECT  353.095 0.17 353.355 12.9 ;
        RECT  353.605 0.17 353.865 12.9 ;
        RECT  352.585 0.52 352.845 5.815 ;
        RECT  353.17 190.585 353.37 191.315 ;
        RECT  354.115 0.17 354.885 0.43 ;
        RECT  354.115 0.17 354.375 11.5 ;
        RECT  354.625 0.17 354.885 11.5 ;
        RECT  353.665 190.585 353.865 191.315 ;
        RECT  354.165 190.585 354.365 191.315 ;
        RECT  354.665 190.585 354.865 191.315 ;
        RECT  356.155 0.17 356.925 0.43 ;
        RECT  356.155 0.17 356.415 10.48 ;
        RECT  356.665 0.17 356.925 10.99 ;
        RECT  355.16 190.585 355.36 191.315 ;
        RECT  355.98 190.585 356.18 191.315 ;
        RECT  357.175 0.17 357.945 0.94 ;
        RECT  357.175 0.17 357.435 8.7 ;
        RECT  357.685 0.17 357.945 12.9 ;
        RECT  356.475 190.585 356.675 191.315 ;
        RECT  356.975 190.585 357.175 191.315 ;
        RECT  357.475 190.585 357.675 191.315 ;
        RECT  357.97 190.585 358.17 191.315 ;
        RECT  358.195 0.52 358.455 2.485 ;
        RECT  358.79 190.585 358.99 191.315 ;
        RECT  359.06 0.52 359.32 14.11 ;
        RECT  359.285 190.585 359.485 191.315 ;
        RECT  359.57 0.52 359.83 2.335 ;
        RECT  359.785 190.585 359.985 191.315 ;
        RECT  360.285 190.585 360.485 191.315 ;
        RECT  362.275 0.17 363.045 0.43 ;
        RECT  362.275 0.17 362.535 8.7 ;
        RECT  362.785 0.17 363.045 8.7 ;
        RECT  363.295 0.17 364.065 0.94 ;
        RECT  363.295 0.17 363.555 8.7 ;
        RECT  363.805 0.17 364.065 8.7 ;
        RECT  364.315 0.17 365.085 0.43 ;
        RECT  364.315 0.17 364.575 8.7 ;
        RECT  364.825 0.17 365.085 8.7 ;
        RECT  365.335 0.17 366.105 0.94 ;
        RECT  365.335 0.17 365.595 8.7 ;
        RECT  365.845 0.17 366.105 8.7 ;
        RECT  366.355 0.17 367.125 0.43 ;
        RECT  366.355 0.17 366.615 8.7 ;
        RECT  366.865 0.17 367.125 8.7 ;
        RECT  367.375 0.17 368.145 0.94 ;
        RECT  367.375 0.17 367.635 8.7 ;
        RECT  367.885 0.17 368.145 8.7 ;
        RECT  368.395 0.17 369.165 0.43 ;
        RECT  368.395 0.17 368.655 8.7 ;
        RECT  368.905 0.17 369.165 8.7 ;
        RECT  369.415 0.17 370.185 0.94 ;
        RECT  369.415 0.17 369.675 8.7 ;
        RECT  369.925 0.17 370.185 8.7 ;
        RECT  370.435 0.17 371.205 0.43 ;
        RECT  370.435 0.17 370.695 8.7 ;
        RECT  370.945 0.17 371.205 8.7 ;
        RECT  371.455 0.17 372.225 0.94 ;
        RECT  371.455 0.17 371.715 8.7 ;
        RECT  371.965 0.17 372.225 8.7 ;
        RECT  360.78 190.585 360.98 191.315 ;
        RECT  361.6 190.585 361.8 191.315 ;
        RECT  362.595 190.585 362.795 191.315 ;
        RECT  374.16 0.17 374.93 0.94 ;
        RECT  374.16 0.17 374.42 8.7 ;
        RECT  374.67 0.17 374.93 8.7 ;
        RECT  372.63 0.3 372.89 8.7 ;
        RECT  373.14 0 373.4 8.7 ;
        RECT  373.65 0 373.91 8.7 ;
        RECT  375.18 0 375.44 8.7 ;
        RECT  375.69 0 375.95 8.7 ;
        RECT  376.2 0.52 376.46 8.7 ;
        RECT  376.71 0.52 376.97 8.7 ;
        RECT  377.22 0.52 377.48 8.7 ;
        RECT  379.26 0.17 380.03 0.94 ;
        RECT  379.26 0.17 379.52 8.7 ;
        RECT  379.77 0.17 380.03 8.7 ;
        RECT  380.28 0.17 381.05 0.43 ;
        RECT  380.28 0.17 380.54 8.7 ;
        RECT  380.79 0.17 381.05 8.7 ;
        RECT  377.73 0.52 377.99 8.7 ;
        RECT  378.24 0 378.5 8.7 ;
        RECT  378.75 0 379.01 8.7 ;
        RECT  381.3 0.3 381.56 8.7 ;
        RECT  381.81 0.3 382.07 8.7 ;
        RECT  383.85 0.17 384.62 0.94 ;
        RECT  383.85 0.17 384.11 8.7 ;
        RECT  384.36 0.17 384.62 8.7 ;
        RECT  382.32 0.3 382.58 8.7 ;
        RECT  382.83 0.3 383.09 8.7 ;
        RECT  383.34 0.3 383.6 8.7 ;
        RECT  384.87 0.52 385.13 8.7 ;
        RECT  385.38 0.52 385.64 8.7 ;
        RECT  385.89 0.3 386.15 8.7 ;
        RECT  386.4 0.52 386.66 8.7 ;
        RECT  386.91 0.52 387.17 8.7 ;
        RECT  387.42 0.3 387.68 8.7 ;
        RECT  387.93 0.52 388.19 8.7 ;
        RECT  388.44 0.52 388.7 8.7 ;
        RECT  388.95 0.52 389.21 8.7 ;
        RECT  389.46 0.52 389.72 8.7 ;
        RECT  389.97 0.52 390.23 8.7 ;
        RECT  390.48 0.3 390.74 8.7 ;
        RECT  390.99 0.52 391.25 8.7 ;
        RECT  391.5 0.52 391.76 8.7 ;
        RECT  392.01 0.3 392.27 8.7 ;
        RECT  394.05 0.17 394.82 0.94 ;
        RECT  394.05 0.17 394.31 8.7 ;
        RECT  394.56 0.17 394.82 8.7 ;
        RECT  392.52 0.52 392.78 8.7 ;
        RECT  393.03 0.52 393.29 8.7 ;
        RECT  393.54 0.3 393.8 8.7 ;
        RECT  395.07 0.52 395.33 8.7 ;
        RECT  395.58 0.52 395.84 8.7 ;
        RECT  396.09 0.52 396.35 8.7 ;
        RECT  396.6 0.52 396.86 8.7 ;
        RECT  397.11 0.52 397.37 8.7 ;
        RECT  397.62 0.52 397.88 8.7 ;
        RECT  398.13 0.52 398.39 8.7 ;
        RECT  400.17 0.17 400.94 0.94 ;
        RECT  400.17 0.17 400.43 8.7 ;
        RECT  400.68 0.17 400.94 8.7 ;
        RECT  398.64 0.52 398.9 8.7 ;
        RECT  399.15 0 399.41 8.7 ;
        RECT  399.66 0 399.92 8.7 ;
        RECT  401.19 0 401.45 8.7 ;
        RECT  403.23 0.17 404 0.43 ;
        RECT  403.23 0.17 403.49 8.7 ;
        RECT  403.74 0.17 404 8.7 ;
        RECT  401.7 0 401.96 8.7 ;
        RECT  402.21 0.3 402.47 8.7 ;
        RECT  402.72 0.3 402.98 8.7 ;
        RECT  404.25 0.3 404.51 8.7 ;
        RECT  404.76 0.3 405.02 8.7 ;
        RECT  405.27 0.3 405.53 8.7 ;
        RECT  405.78 0.3 406.04 8.7 ;
        RECT  406.29 0.52 406.55 8.7 ;
        RECT  406.8 0.52 407.06 8.7 ;
        RECT  408.84 0.17 409.61 0.43 ;
        RECT  408.84 0.17 409.1 8.7 ;
        RECT  409.35 0.17 409.61 8.7 ;
        RECT  409.86 0.17 410.63 0.94 ;
        RECT  409.86 0.17 410.12 25.5 ;
        RECT  410.37 0.17 410.63 33.9 ;
        RECT  410.88 0.17 411.65 0.43 ;
        RECT  410.88 0.17 411.14 8.7 ;
        RECT  411.39 0.17 411.65 8.7 ;
        RECT  412.255 0.17 413.025 0.94 ;
        RECT  412.255 0.17 412.515 8.7 ;
        RECT  412.765 0.17 413.025 8.7 ;
        RECT  413.275 0.17 414.045 0.43 ;
        RECT  413.275 0.17 413.535 8.7 ;
        RECT  413.785 0.17 414.045 8.7 ;
        RECT  414.295 0.17 415.065 0.94 ;
        RECT  414.295 0.17 414.555 8.7 ;
        RECT  414.805 0.17 415.065 8.7 ;
        RECT  415.315 0.17 416.085 0.43 ;
        RECT  415.315 0.17 415.575 8.7 ;
        RECT  415.825 0.17 416.085 8.7 ;
        RECT  416.335 0.17 417.105 0.94 ;
        RECT  416.335 0.17 416.595 8.7 ;
        RECT  416.845 0.17 417.105 8.7 ;
        RECT  417.355 0.17 418.125 0.43 ;
        RECT  417.355 0.17 417.615 8.7 ;
        RECT  417.865 0.17 418.125 8.7 ;
        RECT  418.375 0.17 419.145 0.94 ;
        RECT  418.375 0.17 418.635 8.7 ;
        RECT  418.885 0.17 419.145 8.7 ;
        RECT  419.395 0.17 420.165 0.43 ;
        RECT  419.395 0.17 419.655 8.7 ;
        RECT  419.905 0.17 420.165 8.7 ;
        RECT  420.415 0.17 421.185 0.94 ;
        RECT  420.415 0.17 420.675 8.7 ;
        RECT  420.925 0.17 421.185 8.7 ;
        RECT  407.31 0.3 407.57 8.7 ;
        RECT  421.435 0.17 422.205 0.43 ;
        RECT  421.435 0.17 421.695 8.7 ;
        RECT  421.945 0.17 422.205 8.7 ;
        RECT  407.82 0.3 408.08 8.7 ;
        RECT  408.33 0.52 408.59 8.7 ;
        RECT  421.685 190.585 421.885 191.315 ;
        RECT  422.68 190.585 422.88 191.315 ;
        RECT  423.5 190.585 423.7 191.315 ;
        RECT  423.995 190.585 424.195 191.315 ;
        RECT  424.495 190.585 424.695 191.315 ;
        RECT  424.65 0.52 424.91 2.335 ;
        RECT  424.995 190.585 425.195 191.315 ;
        RECT  425.16 0.52 425.42 14.11 ;
        RECT  425.49 190.585 425.69 191.315 ;
        RECT  426.535 0.17 427.305 0.94 ;
        RECT  427.045 0.17 427.305 8.7 ;
        RECT  426.535 0.17 426.795 12.9 ;
        RECT  426.025 0.52 426.285 2.485 ;
        RECT  426.31 190.585 426.51 191.315 ;
        RECT  427.555 0.17 428.325 0.43 ;
        RECT  428.065 0.17 428.325 10.48 ;
        RECT  427.555 0.17 427.815 10.99 ;
        RECT  426.805 190.585 427.005 191.315 ;
        RECT  427.305 190.585 427.505 191.315 ;
        RECT  427.805 190.585 428.005 191.315 ;
        RECT  428.3 190.585 428.5 191.315 ;
        RECT  429.595 0.17 430.365 0.43 ;
        RECT  429.595 0.17 429.855 11.5 ;
        RECT  430.105 0.17 430.365 11.5 ;
        RECT  429.12 190.585 429.32 191.315 ;
        RECT  429.615 190.585 429.815 191.315 ;
        RECT  430.615 0.17 431.385 0.94 ;
        RECT  430.615 0.17 430.875 12.9 ;
        RECT  431.125 0.17 431.385 12.9 ;
        RECT  430.115 190.585 430.315 191.315 ;
        RECT  430.615 190.585 430.815 191.315 ;
        RECT  431.11 190.585 431.31 191.315 ;
        RECT  431.635 0.52 431.895 5.815 ;
        RECT  432.49 0.52 432.75 5.16 ;
        RECT  432.49 4.9 433.27 5.16 ;
        RECT  433.01 4.9 433.27 6.64 ;
        RECT  431.93 190.585 432.13 191.315 ;
        RECT  432.425 190.585 432.625 191.315 ;
        RECT  432.925 190.585 433.125 191.315 ;
        RECT  433.425 190.585 433.625 191.315 ;
        RECT  433.92 190.585 434.12 191.315 ;
        RECT  434.74 190.585 434.94 191.315 ;
        RECT  435.235 190.585 435.435 191.315 ;
        RECT  435.735 190.585 435.935 191.315 ;
        RECT  435.89 0.52 436.15 2.335 ;
        RECT  436.235 190.585 436.435 191.315 ;
        RECT  436.4 0.52 436.66 14.11 ;
        RECT  436.73 190.585 436.93 191.315 ;
        RECT  437.775 0.17 438.545 0.94 ;
        RECT  438.285 0.17 438.545 8.7 ;
        RECT  437.775 0.17 438.035 12.9 ;
        RECT  437.265 0.52 437.525 2.485 ;
        RECT  437.55 190.585 437.75 191.315 ;
        RECT  438.795 0.17 439.565 0.43 ;
        RECT  439.305 0.17 439.565 10.48 ;
        RECT  438.795 0.17 439.055 10.99 ;
        RECT  438.045 190.585 438.245 191.315 ;
        RECT  438.545 190.585 438.745 191.315 ;
        RECT  439.045 190.585 439.245 191.315 ;
        RECT  439.54 190.585 439.74 191.315 ;
        RECT  440.835 0.17 441.605 0.43 ;
        RECT  440.835 0.17 441.095 11.5 ;
        RECT  441.345 0.17 441.605 11.5 ;
        RECT  440.36 190.585 440.56 191.315 ;
        RECT  440.855 190.585 441.055 191.315 ;
        RECT  441.855 0.17 442.625 0.94 ;
        RECT  441.855 0.17 442.115 12.9 ;
        RECT  442.365 0.17 442.625 12.9 ;
        RECT  441.355 190.585 441.555 191.315 ;
        RECT  441.855 190.585 442.055 191.315 ;
        RECT  442.35 190.585 442.55 191.315 ;
        RECT  442.875 0.52 443.135 5.815 ;
        RECT  443.73 0.52 443.99 5.16 ;
        RECT  443.73 4.9 444.51 5.16 ;
        RECT  444.25 4.9 444.51 6.64 ;
        RECT  443.17 190.585 443.37 191.315 ;
        RECT  443.665 190.585 443.865 191.315 ;
        RECT  444.165 190.585 444.365 191.315 ;
        RECT  444.665 190.585 444.865 191.315 ;
        RECT  445.16 190.585 445.36 191.315 ;
        RECT  445.98 190.585 446.18 191.315 ;
        RECT  446.475 190.585 446.675 191.315 ;
        RECT  446.975 190.585 447.175 191.315 ;
        RECT  447.13 0.52 447.39 2.335 ;
        RECT  447.475 190.585 447.675 191.315 ;
        RECT  447.64 0.52 447.9 14.11 ;
        RECT  447.97 190.585 448.17 191.315 ;
        RECT  449.015 0.17 449.785 0.94 ;
        RECT  449.525 0.17 449.785 8.7 ;
        RECT  449.015 0.17 449.275 12.9 ;
        RECT  448.505 0.52 448.765 2.485 ;
        RECT  448.79 190.585 448.99 191.315 ;
        RECT  450.035 0.17 450.805 0.43 ;
        RECT  450.545 0.17 450.805 10.48 ;
        RECT  450.035 0.17 450.295 10.99 ;
        RECT  449.285 190.585 449.485 191.315 ;
        RECT  449.785 190.585 449.985 191.315 ;
        RECT  450.285 190.585 450.485 191.315 ;
        RECT  450.78 190.585 450.98 191.315 ;
        RECT  452.075 0.17 452.845 0.43 ;
        RECT  452.075 0.17 452.335 11.5 ;
        RECT  452.585 0.17 452.845 11.5 ;
        RECT  451.6 190.585 451.8 191.315 ;
        RECT  452.095 190.585 452.295 191.315 ;
        RECT  453.095 0.17 453.865 0.94 ;
        RECT  453.095 0.17 453.355 12.9 ;
        RECT  453.605 0.17 453.865 12.9 ;
        RECT  452.595 190.585 452.795 191.315 ;
        RECT  453.095 190.585 453.295 191.315 ;
        RECT  453.59 190.585 453.79 191.315 ;
        RECT  454.115 0.52 454.375 5.815 ;
        RECT  454.97 0.52 455.23 5.16 ;
        RECT  454.97 4.9 455.75 5.16 ;
        RECT  455.49 4.9 455.75 6.64 ;
        RECT  454.41 190.585 454.61 191.315 ;
        RECT  454.905 190.585 455.105 191.315 ;
        RECT  455.405 190.585 455.605 191.315 ;
        RECT  455.905 190.585 456.105 191.315 ;
        RECT  456.4 190.585 456.6 191.315 ;
        RECT  457.22 190.585 457.42 191.315 ;
        RECT  457.715 190.585 457.915 191.315 ;
        RECT  458.215 190.585 458.415 191.315 ;
        RECT  458.37 0.52 458.63 2.335 ;
        RECT  458.715 190.585 458.915 191.315 ;
        RECT  458.88 0.52 459.14 14.11 ;
        RECT  459.21 190.585 459.41 191.315 ;
        RECT  460.255 0.17 461.025 0.94 ;
        RECT  460.765 0.17 461.025 8.7 ;
        RECT  460.255 0.17 460.515 12.9 ;
        RECT  459.745 0.52 460.005 2.485 ;
        RECT  460.03 190.585 460.23 191.315 ;
        RECT  461.275 0.17 462.045 0.43 ;
        RECT  461.785 0.17 462.045 10.48 ;
        RECT  461.275 0.17 461.535 10.99 ;
        RECT  460.525 190.585 460.725 191.315 ;
        RECT  461.025 190.585 461.225 191.315 ;
        RECT  461.525 190.585 461.725 191.315 ;
        RECT  462.02 190.585 462.22 191.315 ;
        RECT  463.315 0.17 464.085 0.43 ;
        RECT  463.315 0.17 463.575 11.5 ;
        RECT  463.825 0.17 464.085 11.5 ;
        RECT  462.84 190.585 463.04 191.315 ;
        RECT  463.335 190.585 463.535 191.315 ;
        RECT  464.335 0.17 465.105 0.94 ;
        RECT  464.335 0.17 464.595 12.9 ;
        RECT  464.845 0.17 465.105 12.9 ;
        RECT  463.835 190.585 464.035 191.315 ;
        RECT  464.335 190.585 464.535 191.315 ;
        RECT  464.83 190.585 465.03 191.315 ;
        RECT  465.355 0.52 465.615 5.815 ;
        RECT  466.21 0.52 466.47 5.16 ;
        RECT  466.21 4.9 466.99 5.16 ;
        RECT  466.73 4.9 466.99 6.64 ;
        RECT  465.65 190.585 465.85 191.315 ;
        RECT  466.145 190.585 466.345 191.315 ;
        RECT  466.645 190.585 466.845 191.315 ;
        RECT  467.145 190.585 467.345 191.315 ;
        RECT  467.64 190.585 467.84 191.315 ;
        RECT  468.46 190.585 468.66 191.315 ;
        RECT  468.955 190.585 469.155 191.315 ;
        RECT  469.455 190.585 469.655 191.315 ;
        RECT  469.61 0.52 469.87 2.335 ;
        RECT  469.955 190.585 470.155 191.315 ;
        RECT  470.12 0.52 470.38 14.11 ;
        RECT  470.45 190.585 470.65 191.315 ;
        RECT  471.495 0.17 472.265 0.94 ;
        RECT  472.005 0.17 472.265 8.7 ;
        RECT  471.495 0.17 471.755 12.9 ;
        RECT  470.985 0.52 471.245 2.485 ;
        RECT  471.27 190.585 471.47 191.315 ;
        RECT  472.515 0.17 473.285 0.43 ;
        RECT  473.025 0.17 473.285 10.48 ;
        RECT  472.515 0.17 472.775 10.99 ;
        RECT  471.765 190.585 471.965 191.315 ;
        RECT  472.265 190.585 472.465 191.315 ;
        RECT  472.765 190.585 472.965 191.315 ;
        RECT  473.26 190.585 473.46 191.315 ;
        RECT  474.555 0.17 475.325 0.43 ;
        RECT  474.555 0.17 474.815 11.5 ;
        RECT  475.065 0.17 475.325 11.5 ;
        RECT  474.08 190.585 474.28 191.315 ;
        RECT  474.575 190.585 474.775 191.315 ;
        RECT  475.575 0.17 476.345 0.94 ;
        RECT  475.575 0.17 475.835 12.9 ;
        RECT  476.085 0.17 476.345 12.9 ;
        RECT  475.075 190.585 475.275 191.315 ;
        RECT  475.575 190.585 475.775 191.315 ;
        RECT  476.07 190.585 476.27 191.315 ;
        RECT  476.595 0.52 476.855 5.815 ;
        RECT  477.45 0.52 477.71 5.16 ;
        RECT  477.45 4.9 478.23 5.16 ;
        RECT  477.97 4.9 478.23 6.64 ;
        RECT  476.89 190.585 477.09 191.315 ;
        RECT  477.385 190.585 477.585 191.315 ;
        RECT  477.885 190.585 478.085 191.315 ;
        RECT  478.385 190.585 478.585 191.315 ;
        RECT  478.88 190.585 479.08 191.315 ;
        RECT  479.7 190.585 479.9 191.315 ;
        RECT  480.195 190.585 480.395 191.315 ;
        RECT  480.695 190.585 480.895 191.315 ;
        RECT  480.85 0.52 481.11 2.335 ;
        RECT  481.195 190.585 481.395 191.315 ;
        RECT  481.36 0.52 481.62 14.11 ;
        RECT  481.69 190.585 481.89 191.315 ;
        RECT  482.735 0.17 483.505 0.94 ;
        RECT  483.245 0.17 483.505 8.7 ;
        RECT  482.735 0.17 482.995 12.9 ;
        RECT  482.225 0.52 482.485 2.485 ;
        RECT  482.51 190.585 482.71 191.315 ;
        RECT  483.755 0.17 484.525 0.43 ;
        RECT  484.265 0.17 484.525 10.48 ;
        RECT  483.755 0.17 484.015 10.99 ;
        RECT  483.005 190.585 483.205 191.315 ;
        RECT  483.505 190.585 483.705 191.315 ;
        RECT  484.005 190.585 484.205 191.315 ;
        RECT  484.5 190.585 484.7 191.315 ;
        RECT  485.795 0.17 486.565 0.43 ;
        RECT  485.795 0.17 486.055 11.5 ;
        RECT  486.305 0.17 486.565 11.5 ;
        RECT  485.32 190.585 485.52 191.315 ;
        RECT  485.815 190.585 486.015 191.315 ;
        RECT  486.815 0.17 487.585 0.94 ;
        RECT  486.815 0.17 487.075 12.9 ;
        RECT  487.325 0.17 487.585 12.9 ;
        RECT  486.315 190.585 486.515 191.315 ;
        RECT  486.815 190.585 487.015 191.315 ;
        RECT  487.31 190.585 487.51 191.315 ;
        RECT  487.835 0.52 488.095 5.815 ;
        RECT  488.69 0.52 488.95 5.16 ;
        RECT  488.69 4.9 489.47 5.16 ;
        RECT  489.21 4.9 489.47 6.64 ;
        RECT  488.13 190.585 488.33 191.315 ;
        RECT  488.625 190.585 488.825 191.315 ;
        RECT  489.125 190.585 489.325 191.315 ;
        RECT  489.625 190.585 489.825 191.315 ;
        RECT  490.12 190.585 490.32 191.315 ;
        RECT  490.94 190.585 491.14 191.315 ;
        RECT  491.435 190.585 491.635 191.315 ;
        RECT  491.935 190.585 492.135 191.315 ;
        RECT  492.09 0.52 492.35 2.335 ;
        RECT  492.435 190.585 492.635 191.315 ;
        RECT  492.6 0.52 492.86 14.11 ;
        RECT  492.93 190.585 493.13 191.315 ;
        RECT  493.975 0.17 494.745 0.94 ;
        RECT  494.485 0.17 494.745 8.7 ;
        RECT  493.975 0.17 494.235 12.9 ;
        RECT  493.465 0.52 493.725 2.485 ;
        RECT  493.75 190.585 493.95 191.315 ;
        RECT  494.995 0.17 495.765 0.43 ;
        RECT  495.505 0.17 495.765 10.48 ;
        RECT  494.995 0.17 495.255 10.99 ;
        RECT  494.245 190.585 494.445 191.315 ;
        RECT  494.745 190.585 494.945 191.315 ;
        RECT  495.245 190.585 495.445 191.315 ;
        RECT  495.74 190.585 495.94 191.315 ;
        RECT  497.035 0.17 497.805 0.43 ;
        RECT  497.035 0.17 497.295 11.5 ;
        RECT  497.545 0.17 497.805 11.5 ;
        RECT  496.56 190.585 496.76 191.315 ;
        RECT  497.055 190.585 497.255 191.315 ;
        RECT  498.055 0.17 498.825 0.94 ;
        RECT  498.055 0.17 498.315 12.9 ;
        RECT  498.565 0.17 498.825 12.9 ;
        RECT  497.555 190.585 497.755 191.315 ;
        RECT  498.055 190.585 498.255 191.315 ;
        RECT  498.55 190.585 498.75 191.315 ;
        RECT  499.075 0.52 499.335 5.815 ;
        RECT  499.93 0.52 500.19 5.16 ;
        RECT  499.93 4.9 500.71 5.16 ;
        RECT  500.45 4.9 500.71 6.64 ;
        RECT  499.37 190.585 499.57 191.315 ;
        RECT  499.865 190.585 500.065 191.315 ;
        RECT  500.365 190.585 500.565 191.315 ;
        RECT  500.865 190.585 501.065 191.315 ;
        RECT  501.36 190.585 501.56 191.315 ;
        RECT  502.18 190.585 502.38 191.315 ;
        RECT  502.675 190.585 502.875 191.315 ;
        RECT  503.175 190.585 503.375 191.315 ;
        RECT  503.33 0.52 503.59 2.335 ;
        RECT  503.675 190.585 503.875 191.315 ;
        RECT  503.84 0.52 504.1 14.11 ;
        RECT  504.17 190.585 504.37 191.315 ;
        RECT  505.215 0.17 505.985 0.94 ;
        RECT  505.725 0.17 505.985 8.7 ;
        RECT  505.215 0.17 505.475 12.9 ;
        RECT  504.705 0.52 504.965 2.485 ;
        RECT  504.99 190.585 505.19 191.315 ;
        RECT  506.235 0.17 507.005 0.43 ;
        RECT  506.745 0.17 507.005 10.48 ;
        RECT  506.235 0.17 506.495 10.99 ;
        RECT  505.485 190.585 505.685 191.315 ;
        RECT  505.985 190.585 506.185 191.315 ;
        RECT  506.485 190.585 506.685 191.315 ;
        RECT  506.98 190.585 507.18 191.315 ;
        RECT  508.275 0.17 509.045 0.43 ;
        RECT  508.275 0.17 508.535 11.5 ;
        RECT  508.785 0.17 509.045 11.5 ;
        RECT  507.8 190.585 508 191.315 ;
        RECT  508.295 190.585 508.495 191.315 ;
        RECT  509.295 0.17 510.065 0.94 ;
        RECT  509.295 0.17 509.555 12.9 ;
        RECT  509.805 0.17 510.065 12.9 ;
        RECT  508.795 190.585 508.995 191.315 ;
        RECT  509.295 190.585 509.495 191.315 ;
        RECT  509.79 190.585 509.99 191.315 ;
        RECT  510.315 0.52 510.575 5.815 ;
        RECT  511.17 0.52 511.43 5.16 ;
        RECT  511.17 4.9 511.95 5.16 ;
        RECT  511.69 4.9 511.95 6.64 ;
        RECT  510.61 190.585 510.81 191.315 ;
        RECT  511.105 190.585 511.305 191.315 ;
        RECT  511.605 190.585 511.805 191.315 ;
        RECT  512.105 190.585 512.305 191.315 ;
        RECT  512.6 190.585 512.8 191.315 ;
        RECT  513.42 190.585 513.62 191.315 ;
        RECT  513.915 190.585 514.115 191.315 ;
        RECT  514.415 190.585 514.615 191.315 ;
        RECT  514.57 0.52 514.83 2.335 ;
        RECT  514.915 190.585 515.115 191.315 ;
        RECT  515.08 0.52 515.34 14.11 ;
        RECT  515.41 190.585 515.61 191.315 ;
        RECT  516.455 0.17 517.225 0.94 ;
        RECT  516.965 0.17 517.225 8.7 ;
        RECT  516.455 0.17 516.715 12.9 ;
        RECT  515.945 0.52 516.205 2.485 ;
        RECT  516.23 190.585 516.43 191.315 ;
        RECT  517.475 0.17 518.245 0.43 ;
        RECT  517.985 0.17 518.245 10.48 ;
        RECT  517.475 0.17 517.735 10.99 ;
        RECT  516.725 190.585 516.925 191.315 ;
        RECT  517.225 190.585 517.425 191.315 ;
        RECT  517.725 190.585 517.925 191.315 ;
        RECT  518.22 190.585 518.42 191.315 ;
        RECT  519.515 0.17 520.285 0.43 ;
        RECT  519.515 0.17 519.775 11.5 ;
        RECT  520.025 0.17 520.285 11.5 ;
        RECT  519.04 190.585 519.24 191.315 ;
        RECT  519.535 190.585 519.735 191.315 ;
        RECT  520.535 0.17 521.305 0.94 ;
        RECT  520.535 0.17 520.795 12.9 ;
        RECT  521.045 0.17 521.305 12.9 ;
        RECT  520.035 190.585 520.235 191.315 ;
        RECT  520.535 190.585 520.735 191.315 ;
        RECT  521.03 190.585 521.23 191.315 ;
        RECT  521.555 0.52 521.815 5.815 ;
        RECT  522.41 0.52 522.67 5.16 ;
        RECT  522.41 4.9 523.19 5.16 ;
        RECT  522.93 4.9 523.19 6.64 ;
        RECT  521.85 190.585 522.05 191.315 ;
        RECT  522.345 190.585 522.545 191.315 ;
        RECT  522.845 190.585 523.045 191.315 ;
        RECT  523.345 190.585 523.545 191.315 ;
        RECT  523.84 190.585 524.04 191.315 ;
        RECT  524.66 190.585 524.86 191.315 ;
        RECT  525.155 190.585 525.355 191.315 ;
        RECT  525.655 190.585 525.855 191.315 ;
        RECT  525.81 0.52 526.07 2.335 ;
        RECT  526.155 190.585 526.355 191.315 ;
        RECT  526.32 0.52 526.58 14.11 ;
        RECT  526.65 190.585 526.85 191.315 ;
        RECT  527.695 0.17 528.465 0.94 ;
        RECT  528.205 0.17 528.465 8.7 ;
        RECT  527.695 0.17 527.955 12.9 ;
        RECT  527.185 0.52 527.445 2.485 ;
        RECT  527.47 190.585 527.67 191.315 ;
        RECT  528.715 0.17 529.485 0.43 ;
        RECT  529.225 0.17 529.485 10.48 ;
        RECT  528.715 0.17 528.975 10.99 ;
        RECT  527.965 190.585 528.165 191.315 ;
        RECT  528.465 190.585 528.665 191.315 ;
        RECT  528.965 190.585 529.165 191.315 ;
        RECT  529.46 190.585 529.66 191.315 ;
        RECT  530.755 0.17 531.525 0.43 ;
        RECT  530.755 0.17 531.015 11.5 ;
        RECT  531.265 0.17 531.525 11.5 ;
        RECT  530.28 190.585 530.48 191.315 ;
        RECT  530.775 190.585 530.975 191.315 ;
        RECT  531.775 0.17 532.545 0.94 ;
        RECT  531.775 0.17 532.035 12.9 ;
        RECT  532.285 0.17 532.545 12.9 ;
        RECT  531.275 190.585 531.475 191.315 ;
        RECT  531.775 190.585 531.975 191.315 ;
        RECT  532.27 190.585 532.47 191.315 ;
        RECT  532.795 0.52 533.055 5.815 ;
        RECT  533.65 0.52 533.91 5.16 ;
        RECT  533.65 4.9 534.43 5.16 ;
        RECT  534.17 4.9 534.43 6.64 ;
        RECT  533.09 190.585 533.29 191.315 ;
        RECT  533.585 190.585 533.785 191.315 ;
        RECT  534.085 190.585 534.285 191.315 ;
        RECT  534.585 190.585 534.785 191.315 ;
        RECT  535.08 190.585 535.28 191.315 ;
        RECT  535.9 190.585 536.1 191.315 ;
        RECT  536.395 190.585 536.595 191.315 ;
        RECT  536.895 190.585 537.095 191.315 ;
        RECT  537.05 0.52 537.31 2.335 ;
        RECT  537.395 190.585 537.595 191.315 ;
        RECT  537.56 0.52 537.82 14.11 ;
        RECT  537.89 190.585 538.09 191.315 ;
        RECT  538.935 0.17 539.705 0.94 ;
        RECT  539.445 0.17 539.705 8.7 ;
        RECT  538.935 0.17 539.195 12.9 ;
        RECT  538.425 0.52 538.685 2.485 ;
        RECT  538.71 190.585 538.91 191.315 ;
        RECT  539.955 0.17 540.725 0.43 ;
        RECT  540.465 0.17 540.725 10.48 ;
        RECT  539.955 0.17 540.215 10.99 ;
        RECT  539.205 190.585 539.405 191.315 ;
        RECT  539.705 190.585 539.905 191.315 ;
        RECT  540.205 190.585 540.405 191.315 ;
        RECT  540.7 190.585 540.9 191.315 ;
        RECT  541.995 0.17 542.765 0.43 ;
        RECT  541.995 0.17 542.255 11.5 ;
        RECT  542.505 0.17 542.765 11.5 ;
        RECT  541.52 190.585 541.72 191.315 ;
        RECT  542.015 190.585 542.215 191.315 ;
        RECT  543.015 0.17 543.785 0.94 ;
        RECT  543.015 0.17 543.275 12.9 ;
        RECT  543.525 0.17 543.785 12.9 ;
        RECT  542.515 190.585 542.715 191.315 ;
        RECT  543.015 190.585 543.215 191.315 ;
        RECT  543.51 190.585 543.71 191.315 ;
        RECT  544.035 0.52 544.295 5.815 ;
        RECT  544.89 0.52 545.15 5.16 ;
        RECT  544.89 4.9 545.67 5.16 ;
        RECT  545.41 4.9 545.67 6.64 ;
        RECT  544.33 190.585 544.53 191.315 ;
        RECT  544.825 190.585 545.025 191.315 ;
        RECT  545.325 190.585 545.525 191.315 ;
        RECT  545.825 190.585 546.025 191.315 ;
        RECT  546.32 190.585 546.52 191.315 ;
        RECT  547.14 190.585 547.34 191.315 ;
        RECT  547.635 190.585 547.835 191.315 ;
        RECT  548.135 190.585 548.335 191.315 ;
        RECT  548.29 0.52 548.55 2.335 ;
        RECT  548.635 190.585 548.835 191.315 ;
        RECT  548.8 0.52 549.06 14.11 ;
        RECT  549.13 190.585 549.33 191.315 ;
        RECT  550.175 0.17 550.945 0.94 ;
        RECT  550.685 0.17 550.945 8.7 ;
        RECT  550.175 0.17 550.435 12.9 ;
        RECT  549.665 0.52 549.925 2.485 ;
        RECT  549.95 190.585 550.15 191.315 ;
        RECT  551.195 0.17 551.965 0.43 ;
        RECT  551.705 0.17 551.965 10.48 ;
        RECT  551.195 0.17 551.455 10.99 ;
        RECT  550.445 190.585 550.645 191.315 ;
        RECT  550.945 190.585 551.145 191.315 ;
        RECT  551.445 190.585 551.645 191.315 ;
        RECT  551.94 190.585 552.14 191.315 ;
        RECT  553.235 0.17 554.005 0.43 ;
        RECT  553.235 0.17 553.495 11.5 ;
        RECT  553.745 0.17 554.005 11.5 ;
        RECT  552.76 190.585 552.96 191.315 ;
        RECT  553.255 190.585 553.455 191.315 ;
        RECT  554.255 0.17 555.025 0.94 ;
        RECT  554.255 0.17 554.515 12.9 ;
        RECT  554.765 0.17 555.025 12.9 ;
        RECT  553.755 190.585 553.955 191.315 ;
        RECT  554.255 190.585 554.455 191.315 ;
        RECT  554.75 190.585 554.95 191.315 ;
        RECT  555.275 0.52 555.535 5.815 ;
        RECT  556.13 0.52 556.39 5.16 ;
        RECT  556.13 4.9 556.91 5.16 ;
        RECT  556.65 4.9 556.91 6.64 ;
        RECT  555.57 190.585 555.77 191.315 ;
        RECT  556.065 190.585 556.265 191.315 ;
        RECT  556.565 190.585 556.765 191.315 ;
        RECT  557.065 190.585 557.265 191.315 ;
        RECT  557.56 190.585 557.76 191.315 ;
        RECT  558.38 190.585 558.58 191.315 ;
        RECT  558.875 190.585 559.075 191.315 ;
        RECT  559.375 190.585 559.575 191.315 ;
        RECT  559.53 0.52 559.79 2.335 ;
        RECT  559.875 190.585 560.075 191.315 ;
        RECT  560.04 0.52 560.3 14.11 ;
        RECT  560.37 190.585 560.57 191.315 ;
        RECT  561.415 0.17 562.185 0.94 ;
        RECT  561.925 0.17 562.185 8.7 ;
        RECT  561.415 0.17 561.675 12.9 ;
        RECT  560.905 0.52 561.165 2.485 ;
        RECT  561.19 190.585 561.39 191.315 ;
        RECT  562.435 0.17 563.205 0.43 ;
        RECT  562.945 0.17 563.205 10.48 ;
        RECT  562.435 0.17 562.695 10.99 ;
        RECT  561.685 190.585 561.885 191.315 ;
        RECT  562.185 190.585 562.385 191.315 ;
        RECT  562.685 190.585 562.885 191.315 ;
        RECT  563.18 190.585 563.38 191.315 ;
        RECT  564.475 0.17 565.245 0.43 ;
        RECT  564.475 0.17 564.735 11.5 ;
        RECT  564.985 0.17 565.245 11.5 ;
        RECT  564 190.585 564.2 191.315 ;
        RECT  564.495 190.585 564.695 191.315 ;
        RECT  565.495 0.17 566.265 0.94 ;
        RECT  565.495 0.17 565.755 12.9 ;
        RECT  566.005 0.17 566.265 12.9 ;
        RECT  564.995 190.585 565.195 191.315 ;
        RECT  565.495 190.585 565.695 191.315 ;
        RECT  565.99 190.585 566.19 191.315 ;
        RECT  566.515 0.52 566.775 5.815 ;
        RECT  567.37 0.52 567.63 5.16 ;
        RECT  567.37 4.9 568.15 5.16 ;
        RECT  567.89 4.9 568.15 6.64 ;
        RECT  566.81 190.585 567.01 191.315 ;
        RECT  567.305 190.585 567.505 191.315 ;
        RECT  567.805 190.585 568.005 191.315 ;
        RECT  568.305 190.585 568.505 191.315 ;
        RECT  568.8 190.585 569 191.315 ;
        RECT  569.62 190.585 569.82 191.315 ;
        RECT  570.115 190.585 570.315 191.315 ;
        RECT  570.615 190.585 570.815 191.315 ;
        RECT  570.77 0.52 571.03 2.335 ;
        RECT  571.115 190.585 571.315 191.315 ;
        RECT  571.28 0.52 571.54 14.11 ;
        RECT  571.61 190.585 571.81 191.315 ;
        RECT  572.655 0.17 573.425 0.94 ;
        RECT  573.165 0.17 573.425 8.7 ;
        RECT  572.655 0.17 572.915 12.9 ;
        RECT  572.145 0.52 572.405 2.485 ;
        RECT  572.43 190.585 572.63 191.315 ;
        RECT  573.675 0.17 574.445 0.43 ;
        RECT  574.185 0.17 574.445 10.48 ;
        RECT  573.675 0.17 573.935 10.99 ;
        RECT  572.925 190.585 573.125 191.315 ;
        RECT  573.425 190.585 573.625 191.315 ;
        RECT  573.925 190.585 574.125 191.315 ;
        RECT  574.42 190.585 574.62 191.315 ;
        RECT  575.715 0.17 576.485 0.43 ;
        RECT  575.715 0.17 575.975 11.5 ;
        RECT  576.225 0.17 576.485 11.5 ;
        RECT  575.24 190.585 575.44 191.315 ;
        RECT  575.735 190.585 575.935 191.315 ;
        RECT  576.735 0.17 577.505 0.94 ;
        RECT  576.735 0.17 576.995 12.9 ;
        RECT  577.245 0.17 577.505 12.9 ;
        RECT  576.235 190.585 576.435 191.315 ;
        RECT  576.735 190.585 576.935 191.315 ;
        RECT  577.23 190.585 577.43 191.315 ;
        RECT  577.755 0.52 578.015 5.815 ;
        RECT  578.61 0.52 578.87 5.16 ;
        RECT  578.61 4.9 579.39 5.16 ;
        RECT  579.13 4.9 579.39 6.64 ;
        RECT  578.05 190.585 578.25 191.315 ;
        RECT  578.545 190.585 578.745 191.315 ;
        RECT  579.045 190.585 579.245 191.315 ;
        RECT  579.545 190.585 579.745 191.315 ;
        RECT  580.04 190.585 580.24 191.315 ;
        RECT  580.86 190.585 581.06 191.315 ;
        RECT  581.355 190.585 581.555 191.315 ;
        RECT  581.855 190.585 582.055 191.315 ;
        RECT  582.01 0.52 582.27 2.335 ;
        RECT  582.355 190.585 582.555 191.315 ;
        RECT  582.52 0.52 582.78 14.11 ;
        RECT  582.85 190.585 583.05 191.315 ;
        RECT  583.895 0.17 584.665 0.94 ;
        RECT  584.405 0.17 584.665 8.7 ;
        RECT  583.895 0.17 584.155 12.9 ;
        RECT  583.385 0.52 583.645 2.485 ;
        RECT  583.67 190.585 583.87 191.315 ;
        RECT  584.915 0.17 585.685 0.43 ;
        RECT  585.425 0.17 585.685 10.48 ;
        RECT  584.915 0.17 585.175 10.99 ;
        RECT  584.165 190.585 584.365 191.315 ;
        RECT  584.665 190.585 584.865 191.315 ;
        RECT  585.165 190.585 585.365 191.315 ;
        RECT  585.66 190.585 585.86 191.315 ;
        RECT  586.955 0.17 587.725 0.43 ;
        RECT  586.955 0.17 587.215 11.5 ;
        RECT  587.465 0.17 587.725 11.5 ;
        RECT  586.48 190.585 586.68 191.315 ;
        RECT  586.975 190.585 587.175 191.315 ;
        RECT  587.975 0.17 588.745 0.94 ;
        RECT  587.975 0.17 588.235 12.9 ;
        RECT  588.485 0.17 588.745 12.9 ;
        RECT  587.475 190.585 587.675 191.315 ;
        RECT  587.975 190.585 588.175 191.315 ;
        RECT  588.47 190.585 588.67 191.315 ;
        RECT  588.995 0.52 589.255 5.815 ;
        RECT  589.85 0.52 590.11 5.16 ;
        RECT  589.85 4.9 590.63 5.16 ;
        RECT  590.37 4.9 590.63 6.64 ;
        RECT  589.29 190.585 589.49 191.315 ;
        RECT  589.785 190.585 589.985 191.315 ;
        RECT  590.285 190.585 590.485 191.315 ;
        RECT  590.785 190.585 590.985 191.315 ;
        RECT  591.28 190.585 591.48 191.315 ;
        RECT  592.1 190.585 592.3 191.315 ;
        RECT  592.595 190.585 592.795 191.315 ;
        RECT  593.095 190.585 593.295 191.315 ;
        RECT  593.25 0.52 593.51 2.335 ;
        RECT  593.595 190.585 593.795 191.315 ;
        RECT  593.76 0.52 594.02 14.11 ;
        RECT  594.09 190.585 594.29 191.315 ;
        RECT  595.135 0.17 595.905 0.94 ;
        RECT  595.645 0.17 595.905 8.7 ;
        RECT  595.135 0.17 595.395 12.9 ;
        RECT  594.625 0.52 594.885 2.485 ;
        RECT  594.91 190.585 595.11 191.315 ;
        RECT  596.155 0.17 596.925 0.43 ;
        RECT  596.665 0.17 596.925 10.48 ;
        RECT  596.155 0.17 596.415 10.99 ;
        RECT  595.405 190.585 595.605 191.315 ;
        RECT  595.905 190.585 596.105 191.315 ;
        RECT  596.405 190.585 596.605 191.315 ;
        RECT  596.9 190.585 597.1 191.315 ;
        RECT  598.195 0.17 598.965 0.43 ;
        RECT  598.195 0.17 598.455 11.5 ;
        RECT  598.705 0.17 598.965 11.5 ;
        RECT  597.72 190.585 597.92 191.315 ;
        RECT  598.215 190.585 598.415 191.315 ;
        RECT  599.215 0.17 599.985 0.94 ;
        RECT  599.215 0.17 599.475 12.9 ;
        RECT  599.725 0.17 599.985 12.9 ;
        RECT  598.715 190.585 598.915 191.315 ;
        RECT  599.215 190.585 599.415 191.315 ;
        RECT  599.71 190.585 599.91 191.315 ;
        RECT  600.235 0.52 600.495 5.815 ;
        RECT  601.09 0.52 601.35 5.16 ;
        RECT  601.09 4.9 601.87 5.16 ;
        RECT  601.61 4.9 601.87 6.64 ;
        RECT  600.53 190.585 600.73 191.315 ;
        RECT  601.025 190.585 601.225 191.315 ;
        RECT  601.525 190.585 601.725 191.315 ;
        RECT  602.025 190.585 602.225 191.315 ;
        RECT  602.52 190.585 602.72 191.315 ;
        RECT  603.34 190.585 603.54 191.315 ;
        RECT  603.835 190.585 604.035 191.315 ;
        RECT  604.335 190.585 604.535 191.315 ;
        RECT  604.49 0.52 604.75 2.335 ;
        RECT  604.835 190.585 605.035 191.315 ;
        RECT  605 0.52 605.26 14.11 ;
        RECT  605.33 190.585 605.53 191.315 ;
        RECT  606.375 0.17 607.145 0.94 ;
        RECT  606.885 0.17 607.145 8.7 ;
        RECT  606.375 0.17 606.635 12.9 ;
        RECT  605.865 0.52 606.125 2.485 ;
        RECT  606.15 190.585 606.35 191.315 ;
        RECT  607.395 0.17 608.165 0.43 ;
        RECT  607.905 0.17 608.165 10.48 ;
        RECT  607.395 0.17 607.655 10.99 ;
        RECT  606.645 190.585 606.845 191.315 ;
        RECT  607.145 190.585 607.345 191.315 ;
        RECT  607.645 190.585 607.845 191.315 ;
        RECT  608.14 190.585 608.34 191.315 ;
        RECT  609.435 0.17 610.205 0.43 ;
        RECT  609.435 0.17 609.695 11.5 ;
        RECT  609.945 0.17 610.205 11.5 ;
        RECT  608.96 190.585 609.16 191.315 ;
        RECT  609.455 190.585 609.655 191.315 ;
        RECT  610.455 0.17 611.225 0.94 ;
        RECT  610.455 0.17 610.715 12.9 ;
        RECT  610.965 0.17 611.225 12.9 ;
        RECT  609.955 190.585 610.155 191.315 ;
        RECT  610.455 190.585 610.655 191.315 ;
        RECT  610.95 190.585 611.15 191.315 ;
        RECT  611.475 0.52 611.735 5.815 ;
        RECT  612.33 0.52 612.59 5.16 ;
        RECT  612.33 4.9 613.11 5.16 ;
        RECT  612.85 4.9 613.11 6.64 ;
        RECT  611.77 190.585 611.97 191.315 ;
        RECT  612.265 190.585 612.465 191.315 ;
        RECT  612.765 190.585 612.965 191.315 ;
        RECT  613.265 190.585 613.465 191.315 ;
        RECT  613.76 190.585 613.96 191.315 ;
        RECT  614.58 190.585 614.78 191.315 ;
        RECT  615.075 190.585 615.275 191.315 ;
        RECT  615.575 190.585 615.775 191.315 ;
        RECT  615.73 0.52 615.99 2.335 ;
        RECT  616.075 190.585 616.275 191.315 ;
        RECT  616.24 0.52 616.5 14.11 ;
        RECT  616.57 190.585 616.77 191.315 ;
        RECT  617.615 0.17 618.385 0.94 ;
        RECT  618.125 0.17 618.385 8.7 ;
        RECT  617.615 0.17 617.875 12.9 ;
        RECT  617.105 0.52 617.365 2.485 ;
        RECT  617.39 190.585 617.59 191.315 ;
        RECT  618.635 0.17 619.405 0.43 ;
        RECT  619.145 0.17 619.405 10.48 ;
        RECT  618.635 0.17 618.895 10.99 ;
        RECT  617.885 190.585 618.085 191.315 ;
        RECT  618.385 190.585 618.585 191.315 ;
        RECT  618.885 190.585 619.085 191.315 ;
        RECT  619.38 190.585 619.58 191.315 ;
        RECT  620.675 0.17 621.445 0.43 ;
        RECT  620.675 0.17 620.935 11.5 ;
        RECT  621.185 0.17 621.445 11.5 ;
        RECT  620.2 190.585 620.4 191.315 ;
        RECT  620.695 190.585 620.895 191.315 ;
        RECT  621.695 0.17 622.465 0.94 ;
        RECT  621.695 0.17 621.955 12.9 ;
        RECT  622.205 0.17 622.465 12.9 ;
        RECT  621.195 190.585 621.395 191.315 ;
        RECT  621.695 190.585 621.895 191.315 ;
        RECT  622.19 190.585 622.39 191.315 ;
        RECT  622.715 0.52 622.975 5.815 ;
        RECT  623.57 0.52 623.83 5.16 ;
        RECT  623.57 4.9 624.35 5.16 ;
        RECT  624.09 4.9 624.35 6.64 ;
        RECT  623.01 190.585 623.21 191.315 ;
        RECT  623.505 190.585 623.705 191.315 ;
        RECT  624.005 190.585 624.205 191.315 ;
        RECT  624.505 190.585 624.705 191.315 ;
        RECT  625 190.585 625.2 191.315 ;
        RECT  625.82 190.585 626.02 191.315 ;
        RECT  626.315 190.585 626.515 191.315 ;
        RECT  626.815 190.585 627.015 191.315 ;
        RECT  626.97 0.52 627.23 2.335 ;
        RECT  627.315 190.585 627.515 191.315 ;
        RECT  627.48 0.52 627.74 14.11 ;
        RECT  627.81 190.585 628.01 191.315 ;
        RECT  628.855 0.17 629.625 0.94 ;
        RECT  629.365 0.17 629.625 8.7 ;
        RECT  628.855 0.17 629.115 12.9 ;
        RECT  628.345 0.52 628.605 2.485 ;
        RECT  628.63 190.585 628.83 191.315 ;
        RECT  629.875 0.17 630.645 0.43 ;
        RECT  630.385 0.17 630.645 10.48 ;
        RECT  629.875 0.17 630.135 10.99 ;
        RECT  629.125 190.585 629.325 191.315 ;
        RECT  629.625 190.585 629.825 191.315 ;
        RECT  630.125 190.585 630.325 191.315 ;
        RECT  630.62 190.585 630.82 191.315 ;
        RECT  631.915 0.17 632.685 0.43 ;
        RECT  631.915 0.17 632.175 11.5 ;
        RECT  632.425 0.17 632.685 11.5 ;
        RECT  631.44 190.585 631.64 191.315 ;
        RECT  631.935 190.585 632.135 191.315 ;
        RECT  632.935 0.17 633.705 0.94 ;
        RECT  632.935 0.17 633.195 12.9 ;
        RECT  633.445 0.17 633.705 12.9 ;
        RECT  632.435 190.585 632.635 191.315 ;
        RECT  632.935 190.585 633.135 191.315 ;
        RECT  633.43 190.585 633.63 191.315 ;
        RECT  633.955 0.52 634.215 5.815 ;
        RECT  634.81 0.52 635.07 5.16 ;
        RECT  634.81 4.9 635.59 5.16 ;
        RECT  635.33 4.9 635.59 6.64 ;
        RECT  634.25 190.585 634.45 191.315 ;
        RECT  634.745 190.585 634.945 191.315 ;
        RECT  635.245 190.585 635.445 191.315 ;
        RECT  635.745 190.585 635.945 191.315 ;
        RECT  636.24 190.585 636.44 191.315 ;
        RECT  637.06 190.585 637.26 191.315 ;
        RECT  637.555 190.585 637.755 191.315 ;
        RECT  638.055 190.585 638.255 191.315 ;
        RECT  638.21 0.52 638.47 2.335 ;
        RECT  638.555 190.585 638.755 191.315 ;
        RECT  638.72 0.52 638.98 14.11 ;
        RECT  639.05 190.585 639.25 191.315 ;
        RECT  640.095 0.17 640.865 0.94 ;
        RECT  640.605 0.17 640.865 8.7 ;
        RECT  640.095 0.17 640.355 12.9 ;
        RECT  639.585 0.52 639.845 2.485 ;
        RECT  639.87 190.585 640.07 191.315 ;
        RECT  641.115 0.17 641.885 0.43 ;
        RECT  641.625 0.17 641.885 10.48 ;
        RECT  641.115 0.17 641.375 10.99 ;
        RECT  640.365 190.585 640.565 191.315 ;
        RECT  640.865 190.585 641.065 191.315 ;
        RECT  641.365 190.585 641.565 191.315 ;
        RECT  641.86 190.585 642.06 191.315 ;
        RECT  643.155 0.17 643.925 0.43 ;
        RECT  643.155 0.17 643.415 11.5 ;
        RECT  643.665 0.17 643.925 11.5 ;
        RECT  642.68 190.585 642.88 191.315 ;
        RECT  643.175 190.585 643.375 191.315 ;
        RECT  644.175 0.17 644.945 0.94 ;
        RECT  644.175 0.17 644.435 12.9 ;
        RECT  644.685 0.17 644.945 12.9 ;
        RECT  643.675 190.585 643.875 191.315 ;
        RECT  644.175 190.585 644.375 191.315 ;
        RECT  644.67 190.585 644.87 191.315 ;
        RECT  645.195 0.52 645.455 5.815 ;
        RECT  646.05 0.52 646.31 5.16 ;
        RECT  646.05 4.9 646.83 5.16 ;
        RECT  646.57 4.9 646.83 6.64 ;
        RECT  645.49 190.585 645.69 191.315 ;
        RECT  645.985 190.585 646.185 191.315 ;
        RECT  646.485 190.585 646.685 191.315 ;
        RECT  646.985 190.585 647.185 191.315 ;
        RECT  647.48 190.585 647.68 191.315 ;
        RECT  648.3 190.585 648.5 191.315 ;
        RECT  648.795 190.585 648.995 191.315 ;
        RECT  649.295 190.585 649.495 191.315 ;
        RECT  649.45 0.52 649.71 2.335 ;
        RECT  649.795 190.585 649.995 191.315 ;
        RECT  649.96 0.52 650.22 14.11 ;
        RECT  650.29 190.585 650.49 191.315 ;
        RECT  651.335 0.17 652.105 0.94 ;
        RECT  651.845 0.17 652.105 8.7 ;
        RECT  651.335 0.17 651.595 12.9 ;
        RECT  650.825 0.52 651.085 2.485 ;
        RECT  651.11 190.585 651.31 191.315 ;
        RECT  652.355 0.17 653.125 0.43 ;
        RECT  652.865 0.17 653.125 10.48 ;
        RECT  652.355 0.17 652.615 10.99 ;
        RECT  651.605 190.585 651.805 191.315 ;
        RECT  652.105 190.585 652.305 191.315 ;
        RECT  652.605 190.585 652.805 191.315 ;
        RECT  653.1 190.585 653.3 191.315 ;
        RECT  654.395 0.17 655.165 0.43 ;
        RECT  654.395 0.17 654.655 11.5 ;
        RECT  654.905 0.17 655.165 11.5 ;
        RECT  653.92 190.585 654.12 191.315 ;
        RECT  654.415 190.585 654.615 191.315 ;
        RECT  655.415 0.17 656.185 0.94 ;
        RECT  655.415 0.17 655.675 12.9 ;
        RECT  655.925 0.17 656.185 12.9 ;
        RECT  654.915 190.585 655.115 191.315 ;
        RECT  655.415 190.585 655.615 191.315 ;
        RECT  655.91 190.585 656.11 191.315 ;
        RECT  656.435 0.52 656.695 5.815 ;
        RECT  657.29 0.52 657.55 5.16 ;
        RECT  657.29 4.9 658.07 5.16 ;
        RECT  657.81 4.9 658.07 6.64 ;
        RECT  656.73 190.585 656.93 191.315 ;
        RECT  657.225 190.585 657.425 191.315 ;
        RECT  657.725 190.585 657.925 191.315 ;
        RECT  658.225 190.585 658.425 191.315 ;
        RECT  658.72 190.585 658.92 191.315 ;
        RECT  659.54 190.585 659.74 191.315 ;
        RECT  660.035 190.585 660.235 191.315 ;
        RECT  660.535 190.585 660.735 191.315 ;
        RECT  660.69 0.52 660.95 2.335 ;
        RECT  661.035 190.585 661.235 191.315 ;
        RECT  661.2 0.52 661.46 14.11 ;
        RECT  661.53 190.585 661.73 191.315 ;
        RECT  662.575 0.17 663.345 0.94 ;
        RECT  663.085 0.17 663.345 8.7 ;
        RECT  662.575 0.17 662.835 12.9 ;
        RECT  662.065 0.52 662.325 2.485 ;
        RECT  662.35 190.585 662.55 191.315 ;
        RECT  663.595 0.17 664.365 0.43 ;
        RECT  664.105 0.17 664.365 10.48 ;
        RECT  663.595 0.17 663.855 10.99 ;
        RECT  662.845 190.585 663.045 191.315 ;
        RECT  663.345 190.585 663.545 191.315 ;
        RECT  663.845 190.585 664.045 191.315 ;
        RECT  664.34 190.585 664.54 191.315 ;
        RECT  665.635 0.17 666.405 0.43 ;
        RECT  665.635 0.17 665.895 11.5 ;
        RECT  666.145 0.17 666.405 11.5 ;
        RECT  665.16 190.585 665.36 191.315 ;
        RECT  665.655 190.585 665.855 191.315 ;
        RECT  666.655 0.17 667.425 0.94 ;
        RECT  666.655 0.17 666.915 12.9 ;
        RECT  667.165 0.17 667.425 12.9 ;
        RECT  666.155 190.585 666.355 191.315 ;
        RECT  666.655 190.585 666.855 191.315 ;
        RECT  667.15 190.585 667.35 191.315 ;
        RECT  667.675 0.52 667.935 5.815 ;
        RECT  668.53 0.52 668.79 5.16 ;
        RECT  668.53 4.9 669.31 5.16 ;
        RECT  669.05 4.9 669.31 6.64 ;
        RECT  667.97 190.585 668.17 191.315 ;
        RECT  668.465 190.585 668.665 191.315 ;
        RECT  668.965 190.585 669.165 191.315 ;
        RECT  669.465 190.585 669.665 191.315 ;
        RECT  669.96 190.585 670.16 191.315 ;
        RECT  670.78 190.585 670.98 191.315 ;
        RECT  671.275 190.585 671.475 191.315 ;
        RECT  671.775 190.585 671.975 191.315 ;
        RECT  671.93 0.52 672.19 2.335 ;
        RECT  672.275 190.585 672.475 191.315 ;
        RECT  672.44 0.52 672.7 14.11 ;
        RECT  672.77 190.585 672.97 191.315 ;
        RECT  673.815 0.17 674.585 0.94 ;
        RECT  674.325 0.17 674.585 8.7 ;
        RECT  673.815 0.17 674.075 12.9 ;
        RECT  673.305 0.52 673.565 2.485 ;
        RECT  673.59 190.585 673.79 191.315 ;
        RECT  674.835 0.17 675.605 0.43 ;
        RECT  675.345 0.17 675.605 10.48 ;
        RECT  674.835 0.17 675.095 10.99 ;
        RECT  674.085 190.585 674.285 191.315 ;
        RECT  674.585 190.585 674.785 191.315 ;
        RECT  675.085 190.585 675.285 191.315 ;
        RECT  675.58 190.585 675.78 191.315 ;
        RECT  676.875 0.17 677.645 0.43 ;
        RECT  676.875 0.17 677.135 11.5 ;
        RECT  677.385 0.17 677.645 11.5 ;
        RECT  676.4 190.585 676.6 191.315 ;
        RECT  676.895 190.585 677.095 191.315 ;
        RECT  677.895 0.17 678.665 0.94 ;
        RECT  677.895 0.17 678.155 12.9 ;
        RECT  678.405 0.17 678.665 12.9 ;
        RECT  677.395 190.585 677.595 191.315 ;
        RECT  677.895 190.585 678.095 191.315 ;
        RECT  678.39 190.585 678.59 191.315 ;
        RECT  678.915 0.52 679.175 5.815 ;
        RECT  679.77 0.52 680.03 5.16 ;
        RECT  679.77 4.9 680.55 5.16 ;
        RECT  680.29 4.9 680.55 6.64 ;
        RECT  679.21 190.585 679.41 191.315 ;
        RECT  679.705 190.585 679.905 191.315 ;
        RECT  680.205 190.585 680.405 191.315 ;
        RECT  680.705 190.585 680.905 191.315 ;
        RECT  681.2 190.585 681.4 191.315 ;
        RECT  682.02 190.585 682.22 191.315 ;
        RECT  682.515 190.585 682.715 191.315 ;
        RECT  683.015 190.585 683.215 191.315 ;
        RECT  683.17 0.52 683.43 2.335 ;
        RECT  683.515 190.585 683.715 191.315 ;
        RECT  683.68 0.52 683.94 14.11 ;
        RECT  684.01 190.585 684.21 191.315 ;
        RECT  685.055 0.17 685.825 0.94 ;
        RECT  685.565 0.17 685.825 8.7 ;
        RECT  685.055 0.17 685.315 12.9 ;
        RECT  684.545 0.52 684.805 2.485 ;
        RECT  684.83 190.585 685.03 191.315 ;
        RECT  686.075 0.17 686.845 0.43 ;
        RECT  686.585 0.17 686.845 10.48 ;
        RECT  686.075 0.17 686.335 10.99 ;
        RECT  685.325 190.585 685.525 191.315 ;
        RECT  685.825 190.585 686.025 191.315 ;
        RECT  686.325 190.585 686.525 191.315 ;
        RECT  686.82 190.585 687.02 191.315 ;
        RECT  688.115 0.17 688.885 0.43 ;
        RECT  688.115 0.17 688.375 11.5 ;
        RECT  688.625 0.17 688.885 11.5 ;
        RECT  687.64 190.585 687.84 191.315 ;
        RECT  688.135 190.585 688.335 191.315 ;
        RECT  689.135 0.17 689.905 0.94 ;
        RECT  689.135 0.17 689.395 12.9 ;
        RECT  689.645 0.17 689.905 12.9 ;
        RECT  688.635 190.585 688.835 191.315 ;
        RECT  689.135 190.585 689.335 191.315 ;
        RECT  689.63 190.585 689.83 191.315 ;
        RECT  690.155 0.52 690.415 5.815 ;
        RECT  691.01 0.52 691.27 5.16 ;
        RECT  691.01 4.9 691.79 5.16 ;
        RECT  691.53 4.9 691.79 6.64 ;
        RECT  690.45 190.585 690.65 191.315 ;
        RECT  690.945 190.585 691.145 191.315 ;
        RECT  691.445 190.585 691.645 191.315 ;
        RECT  691.945 190.585 692.145 191.315 ;
        RECT  692.44 190.585 692.64 191.315 ;
        RECT  693.26 190.585 693.46 191.315 ;
        RECT  693.755 190.585 693.955 191.315 ;
        RECT  694.255 190.585 694.455 191.315 ;
        RECT  694.41 0.52 694.67 2.335 ;
        RECT  694.755 190.585 694.955 191.315 ;
        RECT  694.92 0.52 695.18 14.11 ;
        RECT  695.25 190.585 695.45 191.315 ;
        RECT  696.295 0.17 697.065 0.94 ;
        RECT  696.805 0.17 697.065 8.7 ;
        RECT  696.295 0.17 696.555 12.9 ;
        RECT  695.785 0.52 696.045 2.485 ;
        RECT  696.07 190.585 696.27 191.315 ;
        RECT  697.315 0.17 698.085 0.43 ;
        RECT  697.825 0.17 698.085 10.48 ;
        RECT  697.315 0.17 697.575 10.99 ;
        RECT  696.565 190.585 696.765 191.315 ;
        RECT  697.065 190.585 697.265 191.315 ;
        RECT  697.565 190.585 697.765 191.315 ;
        RECT  698.06 190.585 698.26 191.315 ;
        RECT  699.355 0.17 700.125 0.43 ;
        RECT  699.355 0.17 699.615 11.5 ;
        RECT  699.865 0.17 700.125 11.5 ;
        RECT  698.88 190.585 699.08 191.315 ;
        RECT  699.375 190.585 699.575 191.315 ;
        RECT  700.375 0.17 701.145 0.94 ;
        RECT  700.375 0.17 700.635 12.9 ;
        RECT  700.885 0.17 701.145 12.9 ;
        RECT  699.875 190.585 700.075 191.315 ;
        RECT  700.375 190.585 700.575 191.315 ;
        RECT  700.87 190.585 701.07 191.315 ;
        RECT  701.395 0.52 701.655 5.815 ;
        RECT  702.25 0.52 702.51 5.16 ;
        RECT  702.25 4.9 703.03 5.16 ;
        RECT  702.77 4.9 703.03 6.64 ;
        RECT  701.69 190.585 701.89 191.315 ;
        RECT  702.185 190.585 702.385 191.315 ;
        RECT  702.685 190.585 702.885 191.315 ;
        RECT  703.185 190.585 703.385 191.315 ;
        RECT  703.68 190.585 703.88 191.315 ;
        RECT  704.5 190.585 704.7 191.315 ;
        RECT  704.995 190.585 705.195 191.315 ;
        RECT  705.495 190.585 705.695 191.315 ;
        RECT  705.65 0.52 705.91 2.335 ;
        RECT  705.995 190.585 706.195 191.315 ;
        RECT  706.16 0.52 706.42 14.11 ;
        RECT  706.49 190.585 706.69 191.315 ;
        RECT  707.535 0.17 708.305 0.94 ;
        RECT  708.045 0.17 708.305 8.7 ;
        RECT  707.535 0.17 707.795 12.9 ;
        RECT  707.025 0.52 707.285 2.485 ;
        RECT  707.31 190.585 707.51 191.315 ;
        RECT  708.555 0.17 709.325 0.43 ;
        RECT  709.065 0.17 709.325 10.48 ;
        RECT  708.555 0.17 708.815 10.99 ;
        RECT  707.805 190.585 708.005 191.315 ;
        RECT  708.305 190.585 708.505 191.315 ;
        RECT  708.805 190.585 709.005 191.315 ;
        RECT  709.3 190.585 709.5 191.315 ;
        RECT  710.595 0.17 711.365 0.43 ;
        RECT  710.595 0.17 710.855 11.5 ;
        RECT  711.105 0.17 711.365 11.5 ;
        RECT  710.12 190.585 710.32 191.315 ;
        RECT  710.615 190.585 710.815 191.315 ;
        RECT  711.615 0.17 712.385 0.94 ;
        RECT  711.615 0.17 711.875 12.9 ;
        RECT  712.125 0.17 712.385 12.9 ;
        RECT  711.115 190.585 711.315 191.315 ;
        RECT  711.615 190.585 711.815 191.315 ;
        RECT  712.11 190.585 712.31 191.315 ;
        RECT  712.635 0.52 712.895 5.815 ;
        RECT  713.49 0.52 713.75 5.16 ;
        RECT  713.49 4.9 714.27 5.16 ;
        RECT  714.01 4.9 714.27 6.64 ;
        RECT  712.93 190.585 713.13 191.315 ;
        RECT  713.425 190.585 713.625 191.315 ;
        RECT  713.925 190.585 714.125 191.315 ;
        RECT  714.425 190.585 714.625 191.315 ;
        RECT  714.92 190.585 715.12 191.315 ;
        RECT  715.74 190.585 715.94 191.315 ;
        RECT  716.235 190.585 716.435 191.315 ;
        RECT  716.735 190.585 716.935 191.315 ;
        RECT  716.89 0.52 717.15 2.335 ;
        RECT  717.235 190.585 717.435 191.315 ;
        RECT  717.4 0.52 717.66 14.11 ;
        RECT  717.73 190.585 717.93 191.315 ;
        RECT  718.775 0.17 719.545 0.94 ;
        RECT  719.285 0.17 719.545 8.7 ;
        RECT  718.775 0.17 719.035 12.9 ;
        RECT  718.265 0.52 718.525 2.485 ;
        RECT  718.55 190.585 718.75 191.315 ;
        RECT  719.795 0.17 720.565 0.43 ;
        RECT  720.305 0.17 720.565 10.48 ;
        RECT  719.795 0.17 720.055 10.99 ;
        RECT  719.045 190.585 719.245 191.315 ;
        RECT  719.545 190.585 719.745 191.315 ;
        RECT  720.045 190.585 720.245 191.315 ;
        RECT  720.54 190.585 720.74 191.315 ;
        RECT  721.835 0.17 722.605 0.43 ;
        RECT  721.835 0.17 722.095 11.5 ;
        RECT  722.345 0.17 722.605 11.5 ;
        RECT  721.36 190.585 721.56 191.315 ;
        RECT  721.855 190.585 722.055 191.315 ;
        RECT  722.855 0.17 723.625 0.94 ;
        RECT  722.855 0.17 723.115 12.9 ;
        RECT  723.365 0.17 723.625 12.9 ;
        RECT  722.355 190.585 722.555 191.315 ;
        RECT  722.855 190.585 723.055 191.315 ;
        RECT  723.35 190.585 723.55 191.315 ;
        RECT  723.875 0.52 724.135 5.815 ;
        RECT  724.73 0.52 724.99 5.16 ;
        RECT  724.73 4.9 725.51 5.16 ;
        RECT  725.25 4.9 725.51 6.64 ;
        RECT  724.17 190.585 724.37 191.315 ;
        RECT  724.665 190.585 724.865 191.315 ;
        RECT  725.165 190.585 725.365 191.315 ;
        RECT  725.665 190.585 725.865 191.315 ;
        RECT  726.16 190.585 726.36 191.315 ;
        RECT  726.98 190.585 727.18 191.315 ;
        RECT  727.475 190.585 727.675 191.315 ;
        RECT  727.975 190.585 728.175 191.315 ;
        RECT  728.13 0.52 728.39 2.335 ;
        RECT  728.475 190.585 728.675 191.315 ;
        RECT  728.64 0.52 728.9 14.11 ;
        RECT  728.97 190.585 729.17 191.315 ;
        RECT  730.015 0.17 730.785 0.94 ;
        RECT  730.525 0.17 730.785 8.7 ;
        RECT  730.015 0.17 730.275 12.9 ;
        RECT  729.505 0.52 729.765 2.485 ;
        RECT  729.79 190.585 729.99 191.315 ;
        RECT  731.035 0.17 731.805 0.43 ;
        RECT  731.545 0.17 731.805 10.48 ;
        RECT  731.035 0.17 731.295 10.99 ;
        RECT  730.285 190.585 730.485 191.315 ;
        RECT  730.785 190.585 730.985 191.315 ;
        RECT  731.285 190.585 731.485 191.315 ;
        RECT  731.78 190.585 731.98 191.315 ;
        RECT  733.075 0.17 733.845 0.43 ;
        RECT  733.075 0.17 733.335 11.5 ;
        RECT  733.585 0.17 733.845 11.5 ;
        RECT  732.6 190.585 732.8 191.315 ;
        RECT  733.095 190.585 733.295 191.315 ;
        RECT  734.095 0.17 734.865 0.94 ;
        RECT  734.095 0.17 734.355 12.9 ;
        RECT  734.605 0.17 734.865 12.9 ;
        RECT  733.595 190.585 733.795 191.315 ;
        RECT  734.095 190.585 734.295 191.315 ;
        RECT  734.59 190.585 734.79 191.315 ;
        RECT  735.115 0.52 735.375 5.815 ;
        RECT  735.97 0.52 736.23 5.16 ;
        RECT  735.97 4.9 736.75 5.16 ;
        RECT  736.49 4.9 736.75 6.64 ;
        RECT  735.41 190.585 735.61 191.315 ;
        RECT  735.905 190.585 736.105 191.315 ;
        RECT  736.405 190.585 736.605 191.315 ;
        RECT  736.905 190.585 737.105 191.315 ;
        RECT  737.4 190.585 737.6 191.315 ;
        RECT  738.22 190.585 738.42 191.315 ;
        RECT  738.715 190.585 738.915 191.315 ;
        RECT  739.215 190.585 739.415 191.315 ;
        RECT  739.37 0.52 739.63 2.335 ;
        RECT  739.715 190.585 739.915 191.315 ;
        RECT  739.88 0.52 740.14 14.11 ;
        RECT  740.21 190.585 740.41 191.315 ;
        RECT  741.255 0.17 742.025 0.94 ;
        RECT  741.765 0.17 742.025 8.7 ;
        RECT  741.255 0.17 741.515 12.9 ;
        RECT  740.745 0.52 741.005 2.485 ;
        RECT  741.03 190.585 741.23 191.315 ;
        RECT  742.275 0.17 743.045 0.43 ;
        RECT  742.785 0.17 743.045 10.48 ;
        RECT  742.275 0.17 742.535 10.99 ;
        RECT  741.525 190.585 741.725 191.315 ;
        RECT  742.025 190.585 742.225 191.315 ;
        RECT  742.525 190.585 742.725 191.315 ;
        RECT  743.02 190.585 743.22 191.315 ;
        RECT  744.315 0.17 745.085 0.43 ;
        RECT  744.315 0.17 744.575 11.5 ;
        RECT  744.825 0.17 745.085 11.5 ;
        RECT  743.84 190.585 744.04 191.315 ;
        RECT  744.335 190.585 744.535 191.315 ;
        RECT  745.335 0.17 746.105 0.94 ;
        RECT  745.335 0.17 745.595 12.9 ;
        RECT  745.845 0.17 746.105 12.9 ;
        RECT  744.835 190.585 745.035 191.315 ;
        RECT  745.335 190.585 745.535 191.315 ;
        RECT  745.83 190.585 746.03 191.315 ;
        RECT  746.355 0.52 746.615 5.815 ;
        RECT  747.21 0.52 747.47 5.16 ;
        RECT  747.21 4.9 747.99 5.16 ;
        RECT  747.73 4.9 747.99 6.64 ;
        RECT  746.65 190.585 746.85 191.315 ;
        RECT  747.145 190.585 747.345 191.315 ;
        RECT  747.645 190.585 747.845 191.315 ;
        RECT  748.145 190.585 748.345 191.315 ;
        RECT  748.64 190.585 748.84 191.315 ;
        RECT  749.46 190.585 749.66 191.315 ;
        RECT  749.955 190.585 750.155 191.315 ;
        RECT  750.455 190.585 750.655 191.315 ;
        RECT  750.61 0.52 750.87 2.335 ;
        RECT  750.955 190.585 751.155 191.315 ;
        RECT  751.12 0.52 751.38 14.11 ;
        RECT  751.45 190.585 751.65 191.315 ;
        RECT  752.495 0.17 753.265 0.94 ;
        RECT  753.005 0.17 753.265 8.7 ;
        RECT  752.495 0.17 752.755 12.9 ;
        RECT  751.985 0.52 752.245 2.485 ;
        RECT  752.27 190.585 752.47 191.315 ;
        RECT  753.515 0.17 754.285 0.43 ;
        RECT  754.025 0.17 754.285 10.48 ;
        RECT  753.515 0.17 753.775 10.99 ;
        RECT  752.765 190.585 752.965 191.315 ;
        RECT  753.265 190.585 753.465 191.315 ;
        RECT  753.765 190.585 753.965 191.315 ;
        RECT  754.26 190.585 754.46 191.315 ;
        RECT  755.555 0.17 756.325 0.43 ;
        RECT  755.555 0.17 755.815 11.5 ;
        RECT  756.065 0.17 756.325 11.5 ;
        RECT  755.08 190.585 755.28 191.315 ;
        RECT  755.575 190.585 755.775 191.315 ;
        RECT  756.575 0.17 757.345 0.94 ;
        RECT  756.575 0.17 756.835 12.9 ;
        RECT  757.085 0.17 757.345 12.9 ;
        RECT  756.075 190.585 756.275 191.315 ;
        RECT  756.575 190.585 756.775 191.315 ;
        RECT  757.07 190.585 757.27 191.315 ;
        RECT  757.595 0.52 757.855 5.815 ;
        RECT  758.45 0.52 758.71 5.16 ;
        RECT  758.45 4.9 759.23 5.16 ;
        RECT  758.97 4.9 759.23 6.64 ;
        RECT  757.89 190.585 758.09 191.315 ;
        RECT  758.385 190.585 758.585 191.315 ;
        RECT  758.885 190.585 759.085 191.315 ;
        RECT  759.385 190.585 759.585 191.315 ;
        RECT  759.88 190.585 760.08 191.315 ;
        RECT  760.7 190.585 760.9 191.315 ;
        RECT  761.195 190.585 761.395 191.315 ;
        RECT  761.695 190.585 761.895 191.315 ;
        RECT  761.85 0.52 762.11 2.335 ;
        RECT  762.195 190.585 762.395 191.315 ;
        RECT  762.36 0.52 762.62 14.11 ;
        RECT  762.69 190.585 762.89 191.315 ;
        RECT  763.735 0.17 764.505 0.94 ;
        RECT  764.245 0.17 764.505 8.7 ;
        RECT  763.735 0.17 763.995 12.9 ;
        RECT  763.225 0.52 763.485 2.485 ;
        RECT  763.51 190.585 763.71 191.315 ;
        RECT  764.755 0.17 765.525 0.43 ;
        RECT  765.265 0.17 765.525 10.48 ;
        RECT  764.755 0.17 765.015 10.99 ;
        RECT  764.005 190.585 764.205 191.315 ;
        RECT  764.505 190.585 764.705 191.315 ;
        RECT  765.005 190.585 765.205 191.315 ;
        RECT  765.5 190.585 765.7 191.315 ;
        RECT  766.795 0.17 767.565 0.43 ;
        RECT  766.795 0.17 767.055 11.5 ;
        RECT  767.305 0.17 767.565 11.5 ;
        RECT  766.32 190.585 766.52 191.315 ;
        RECT  766.815 190.585 767.015 191.315 ;
        RECT  767.815 0.17 768.585 0.94 ;
        RECT  767.815 0.17 768.075 12.9 ;
        RECT  768.325 0.17 768.585 12.9 ;
        RECT  767.315 190.585 767.515 191.315 ;
        RECT  767.815 190.585 768.015 191.315 ;
        RECT  768.31 190.585 768.51 191.315 ;
        RECT  768.835 0.52 769.095 5.815 ;
        RECT  769.69 0.52 769.95 5.16 ;
        RECT  769.69 4.9 770.47 5.16 ;
        RECT  770.21 4.9 770.47 6.64 ;
        RECT  769.13 190.585 769.33 191.315 ;
        RECT  769.625 190.585 769.825 191.315 ;
        RECT  770.125 190.585 770.325 191.315 ;
        RECT  770.625 190.585 770.825 191.315 ;
        RECT  771.12 190.585 771.32 191.315 ;
        RECT  771.94 190.585 772.14 191.315 ;
        RECT  772.435 190.585 772.635 191.315 ;
        RECT  772.935 190.585 773.135 191.315 ;
        RECT  773.09 0.52 773.35 2.335 ;
        RECT  773.435 190.585 773.635 191.315 ;
        RECT  773.6 0.52 773.86 14.11 ;
        RECT  773.93 190.585 774.13 191.315 ;
        RECT  774.975 0.17 775.745 0.94 ;
        RECT  775.485 0.17 775.745 8.7 ;
        RECT  774.975 0.17 775.235 12.9 ;
        RECT  774.465 0.52 774.725 2.485 ;
        RECT  774.75 190.585 774.95 191.315 ;
        RECT  775.995 0.17 776.765 0.43 ;
        RECT  776.505 0.17 776.765 10.48 ;
        RECT  775.995 0.17 776.255 10.99 ;
        RECT  775.245 190.585 775.445 191.315 ;
        RECT  775.745 190.585 775.945 191.315 ;
        RECT  776.245 190.585 776.445 191.315 ;
        RECT  776.74 190.585 776.94 191.315 ;
        RECT  778.035 0.17 778.805 0.43 ;
        RECT  778.035 0.17 778.295 11.5 ;
        RECT  778.545 0.17 778.805 11.5 ;
        RECT  777.56 190.585 777.76 191.315 ;
        RECT  778.055 190.585 778.255 191.315 ;
        RECT  779.055 0.17 779.825 0.94 ;
        RECT  779.055 0.17 779.315 12.9 ;
        RECT  779.565 0.17 779.825 12.9 ;
        RECT  778.555 190.585 778.755 191.315 ;
        RECT  779.055 190.585 779.255 191.315 ;
        RECT  779.55 190.585 779.75 191.315 ;
        RECT  780.075 0.52 780.335 5.815 ;
        RECT  780.93 0.52 781.19 5.16 ;
        RECT  780.93 4.9 781.71 5.16 ;
        RECT  781.45 4.9 781.71 6.64 ;
        RECT  780.37 190.585 780.57 191.315 ;
        RECT  780.865 190.585 781.065 191.315 ;
        RECT  781.365 190.585 781.565 191.315 ;
        RECT  781.865 190.585 782.065 191.315 ;
        RECT  782.36 190.585 782.56 191.315 ;
        RECT  783.18 190.585 783.38 191.315 ;
        RECT  784.175 45.465 784.375 191.315 ;
        RECT  218.225 0 223.055 191.34 ;
        RECT  229.465 0 234.295 191.34 ;
        RECT  240.705 0 245.535 191.34 ;
        RECT  251.945 0 256.775 191.34 ;
        RECT  263.185 0 268.015 191.34 ;
        RECT  274.425 0 279.255 191.34 ;
        RECT  285.665 0 290.495 191.34 ;
        RECT  296.905 0 301.735 191.34 ;
        RECT  308.145 0 312.975 191.34 ;
        RECT  319.385 0 324.215 191.34 ;
        RECT  330.625 0 335.455 191.34 ;
        RECT  341.865 0 346.695 191.34 ;
        RECT  353.105 0 357.935 191.34 ;
        RECT  378.24 0 384.61 191.34 ;
        RECT  393.55 0 394.81 191.34 ;
        RECT  426.545 0 431.375 191.34 ;
        RECT  437.785 0 442.615 191.34 ;
        RECT  449.025 0 453.855 191.34 ;
        RECT  460.265 0 465.095 191.34 ;
        RECT  471.505 0 476.335 191.34 ;
        RECT  482.745 0 487.575 191.34 ;
        RECT  493.985 0 498.815 191.34 ;
        RECT  505.225 0 510.055 191.34 ;
        RECT  516.465 0 521.295 191.34 ;
        RECT  527.705 0 532.535 191.34 ;
        RECT  538.945 0 543.775 191.34 ;
        RECT  550.185 0 555.015 191.34 ;
        RECT  561.425 0 566.255 191.34 ;
        RECT  572.665 0 577.495 191.34 ;
        RECT  583.905 0 588.735 191.34 ;
        RECT  595.145 0 599.975 191.34 ;
        RECT  606.385 0 611.215 191.34 ;
        RECT  617.625 0 622.455 191.34 ;
        RECT  628.865 0 633.695 191.34 ;
        RECT  640.105 0 644.935 191.34 ;
        RECT  651.345 0 656.175 191.34 ;
        RECT  662.585 0 667.415 191.34 ;
        RECT  673.825 0 678.655 191.34 ;
        RECT  685.065 0 689.895 191.34 ;
        RECT  696.305 0 701.135 191.34 ;
        RECT  707.545 0 712.375 191.34 ;
        RECT  718.785 0 723.615 191.34 ;
        RECT  730.025 0 734.855 191.34 ;
        RECT  741.265 0 746.095 191.34 ;
        RECT  752.505 0 757.335 191.34 ;
        RECT  763.745 0 768.575 191.34 ;
        RECT  774.985 0 779.815 191.34 ;
        RECT  385.9 0 386.14 191.34 ;
        RECT  387.43 0 387.67 191.34 ;
        RECT  390.49 0 390.73 191.34 ;
        RECT  392.02 0 392.26 191.34 ;
        RECT  399.15 0 406.03 191.34 ;
        RECT  407.32 0 408.07 191.34 ;
        RECT  0 0 3.03 191.34 ;
        RECT  4.655 0.17 9.505 191.34 ;
        RECT  11.65 0 14.27 191.34 ;
        RECT  15.895 0.17 20.745 191.34 ;
        RECT  22.89 0 25.51 191.34 ;
        RECT  27.135 0.17 31.985 191.34 ;
        RECT  34.13 0 36.75 191.34 ;
        RECT  38.375 0.17 43.225 191.34 ;
        RECT  45.37 0 47.99 191.34 ;
        RECT  49.615 0.17 54.465 191.34 ;
        RECT  56.61 0 59.23 191.34 ;
        RECT  60.855 0.17 65.705 191.34 ;
        RECT  67.85 0 70.47 191.34 ;
        RECT  72.095 0.17 76.945 191.34 ;
        RECT  79.09 0 81.71 191.34 ;
        RECT  83.335 0.17 88.185 191.34 ;
        RECT  90.33 0 92.95 191.34 ;
        RECT  94.575 0.17 99.425 191.34 ;
        RECT  101.57 0 104.19 191.34 ;
        RECT  105.815 0.17 110.665 191.34 ;
        RECT  112.81 0 115.43 191.34 ;
        RECT  117.055 0.17 121.905 191.34 ;
        RECT  124.05 0 126.67 191.34 ;
        RECT  128.295 0.17 133.145 191.34 ;
        RECT  135.29 0 137.91 191.34 ;
        RECT  139.535 0.17 144.385 191.34 ;
        RECT  146.53 0 149.15 191.34 ;
        RECT  150.775 0.17 155.625 191.34 ;
        RECT  157.77 0 160.39 191.34 ;
        RECT  162.015 0.17 166.865 191.34 ;
        RECT  169.01 0 171.63 191.34 ;
        RECT  173.255 0.17 178.105 191.34 ;
        RECT  180.25 0 182.87 191.34 ;
        RECT  184.495 0.17 189.345 191.34 ;
        RECT  191.49 0 194.11 191.34 ;
        RECT  195.735 0.17 200.585 191.34 ;
        RECT  202.73 0 205.35 191.34 ;
        RECT  206.975 0.17 211.825 191.34 ;
        RECT  213.97 0 216.59 191.34 ;
        RECT  218.215 0.17 223.065 191.34 ;
        RECT  225.21 0 227.83 191.34 ;
        RECT  229.455 0.17 234.305 191.34 ;
        RECT  236.45 0 239.07 191.34 ;
        RECT  240.695 0.17 245.545 191.34 ;
        RECT  247.69 0 250.31 191.34 ;
        RECT  251.935 0.17 256.785 191.34 ;
        RECT  258.93 0 261.55 191.34 ;
        RECT  263.175 0.17 268.025 191.34 ;
        RECT  270.17 0 272.79 191.34 ;
        RECT  274.415 0.17 279.265 191.34 ;
        RECT  281.41 0 284.03 191.34 ;
        RECT  285.655 0.17 290.505 191.34 ;
        RECT  292.65 0 295.27 191.34 ;
        RECT  296.895 0.17 301.745 191.34 ;
        RECT  303.89 0 306.51 191.34 ;
        RECT  308.135 0.17 312.985 191.34 ;
        RECT  315.13 0 317.75 191.34 ;
        RECT  319.375 0.17 324.225 191.34 ;
        RECT  326.37 0 328.99 191.34 ;
        RECT  330.615 0.17 335.465 191.34 ;
        RECT  337.61 0 340.23 191.34 ;
        RECT  341.855 0.17 346.705 191.34 ;
        RECT  348.85 0 351.47 191.34 ;
        RECT  353.095 0.17 357.945 191.34 ;
        RECT  360.09 0 375.95 191.34 ;
        RECT  378.24 0.17 384.62 191.34 ;
        RECT  385.89 0.3 386.15 191.34 ;
        RECT  387.42 0.3 387.68 191.34 ;
        RECT  390.48 0.3 390.74 191.34 ;
        RECT  392.01 0.3 392.27 191.34 ;
        RECT  393.55 0.17 394.82 191.34 ;
        RECT  393.54 0.3 394.82 191.34 ;
        RECT  399.15 0.3 406.04 191.34 ;
        RECT  407.31 0.3 408.08 191.34 ;
        RECT  408.85 0 424.39 191.34 ;
        RECT  408.84 0.17 424.39 191.34 ;
        RECT  426.535 0.17 431.385 191.34 ;
        RECT  433.01 0 435.63 191.34 ;
        RECT  437.775 0.17 442.625 191.34 ;
        RECT  444.25 0 446.87 191.34 ;
        RECT  449.015 0.17 453.865 191.34 ;
        RECT  455.49 0 458.11 191.34 ;
        RECT  460.255 0.17 465.105 191.34 ;
        RECT  466.73 0 469.35 191.34 ;
        RECT  471.495 0.17 476.345 191.34 ;
        RECT  477.97 0 480.59 191.34 ;
        RECT  482.735 0.17 487.585 191.34 ;
        RECT  489.21 0 491.83 191.34 ;
        RECT  493.975 0.17 498.825 191.34 ;
        RECT  500.45 0 503.07 191.34 ;
        RECT  505.215 0.17 510.065 191.34 ;
        RECT  511.69 0 514.31 191.34 ;
        RECT  516.455 0.17 521.305 191.34 ;
        RECT  522.93 0 525.55 191.34 ;
        RECT  527.695 0.17 532.545 191.34 ;
        RECT  534.17 0 536.79 191.34 ;
        RECT  538.935 0.17 543.785 191.34 ;
        RECT  545.41 0 548.03 191.34 ;
        RECT  550.175 0.17 555.025 191.34 ;
        RECT  556.65 0 559.27 191.34 ;
        RECT  561.415 0.17 566.265 191.34 ;
        RECT  567.89 0 570.51 191.34 ;
        RECT  572.655 0.17 577.505 191.34 ;
        RECT  579.13 0 581.75 191.34 ;
        RECT  583.895 0.17 588.745 191.34 ;
        RECT  590.37 0 592.99 191.34 ;
        RECT  595.135 0.17 599.985 191.34 ;
        RECT  601.61 0 604.23 191.34 ;
        RECT  606.375 0.17 611.225 191.34 ;
        RECT  612.85 0 615.47 191.34 ;
        RECT  617.615 0.17 622.465 191.34 ;
        RECT  624.09 0 626.71 191.34 ;
        RECT  628.855 0.17 633.705 191.34 ;
        RECT  635.33 0 637.95 191.34 ;
        RECT  640.095 0.17 644.945 191.34 ;
        RECT  646.57 0 649.19 191.34 ;
        RECT  651.335 0.17 656.185 191.34 ;
        RECT  657.81 0 660.43 191.34 ;
        RECT  662.575 0.17 667.425 191.34 ;
        RECT  669.05 0 671.67 191.34 ;
        RECT  673.815 0.17 678.665 191.34 ;
        RECT  680.29 0 682.91 191.34 ;
        RECT  685.055 0.17 689.905 191.34 ;
        RECT  691.53 0 694.15 191.34 ;
        RECT  696.295 0.17 701.145 191.34 ;
        RECT  702.77 0 705.39 191.34 ;
        RECT  707.535 0.17 712.385 191.34 ;
        RECT  714.01 0 716.63 191.34 ;
        RECT  718.775 0.17 723.625 191.34 ;
        RECT  725.25 0 727.87 191.34 ;
        RECT  730.015 0.17 734.865 191.34 ;
        RECT  736.49 0 739.11 191.34 ;
        RECT  741.255 0.17 746.105 191.34 ;
        RECT  747.73 0 750.35 191.34 ;
        RECT  752.495 0.17 757.345 191.34 ;
        RECT  758.97 0 761.59 191.34 ;
        RECT  763.735 0.17 768.585 191.34 ;
        RECT  770.21 0 772.83 191.34 ;
        RECT  774.975 0.17 779.825 191.34 ;
        RECT  781.45 0 784.48 191.34 ;
        RECT  0 0.52 784.48 191.34 ;
        RECT  4.665 0 9.495 191.34 ;
        RECT  15.905 0 20.735 191.34 ;
        RECT  27.145 0 31.975 191.34 ;
        RECT  38.385 0 43.215 191.34 ;
        RECT  49.625 0 54.455 191.34 ;
        RECT  60.865 0 65.695 191.34 ;
        RECT  72.105 0 76.935 191.34 ;
        RECT  83.345 0 88.175 191.34 ;
        RECT  94.585 0 99.415 191.34 ;
        RECT  105.825 0 110.655 191.34 ;
        RECT  117.065 0 121.895 191.34 ;
        RECT  128.305 0 133.135 191.34 ;
        RECT  139.545 0 144.375 191.34 ;
        RECT  150.785 0 155.615 191.34 ;
        RECT  162.025 0 166.855 191.34 ;
        RECT  173.265 0 178.095 191.34 ;
        RECT  184.505 0 189.335 191.34 ;
        RECT  195.745 0 200.575 191.34 ;
        RECT  206.985 0 211.815 191.34 ;
      LAYER Metal3 ;
        RECT  0 0 784.48 191.34 ;
      LAYER Metal4 ;
        RECT  0 39.085 9.62 45.205 ;
        RECT  0 0 4 191.34 ;
        RECT  7.33 0 9.62 191.34 ;
        RECT  12.95 39.085 20.86 45.205 ;
        RECT  12.95 0 15.24 191.34 ;
        RECT  18.57 0 20.86 191.34 ;
        RECT  24.19 39.085 32.1 45.205 ;
        RECT  24.19 0 26.48 191.34 ;
        RECT  29.81 0 32.1 191.34 ;
        RECT  35.43 39.085 43.34 45.205 ;
        RECT  35.43 0 37.72 191.34 ;
        RECT  41.05 0 43.34 191.34 ;
        RECT  46.67 39.085 54.58 45.205 ;
        RECT  46.67 0 48.96 191.34 ;
        RECT  52.29 0 54.58 191.34 ;
        RECT  57.91 39.085 65.82 45.205 ;
        RECT  57.91 0 60.2 191.34 ;
        RECT  63.53 0 65.82 191.34 ;
        RECT  69.15 39.085 77.06 45.205 ;
        RECT  69.15 0 71.44 191.34 ;
        RECT  74.77 0 77.06 191.34 ;
        RECT  80.39 39.085 88.3 45.205 ;
        RECT  80.39 0 82.68 191.34 ;
        RECT  86.01 0 88.3 191.34 ;
        RECT  91.63 39.085 99.54 45.205 ;
        RECT  91.63 0 93.92 191.34 ;
        RECT  97.25 0 99.54 191.34 ;
        RECT  102.87 39.085 110.78 45.205 ;
        RECT  102.87 0 105.16 191.34 ;
        RECT  108.49 0 110.78 191.34 ;
        RECT  114.11 39.085 122.02 45.205 ;
        RECT  114.11 0 116.4 191.34 ;
        RECT  119.73 0 122.02 191.34 ;
        RECT  125.35 39.085 133.26 45.205 ;
        RECT  125.35 0 127.64 191.34 ;
        RECT  130.97 0 133.26 191.34 ;
        RECT  136.59 39.085 144.5 45.205 ;
        RECT  136.59 0 138.88 191.34 ;
        RECT  142.21 0 144.5 191.34 ;
        RECT  147.83 39.085 155.74 45.205 ;
        RECT  147.83 0 150.12 191.34 ;
        RECT  153.45 0 155.74 191.34 ;
        RECT  159.07 39.085 166.98 45.205 ;
        RECT  159.07 0 161.36 191.34 ;
        RECT  164.69 0 166.98 191.34 ;
        RECT  170.31 39.085 178.22 45.205 ;
        RECT  170.31 0 172.6 191.34 ;
        RECT  175.93 0 178.22 191.34 ;
        RECT  181.55 39.085 189.46 45.205 ;
        RECT  181.55 0 183.84 191.34 ;
        RECT  187.17 0 189.46 191.34 ;
        RECT  192.79 39.085 200.7 45.205 ;
        RECT  192.79 0 195.08 191.34 ;
        RECT  198.41 0 200.7 191.34 ;
        RECT  204.03 39.085 211.94 45.205 ;
        RECT  204.03 0 206.32 191.34 ;
        RECT  209.65 0 211.94 191.34 ;
        RECT  215.27 39.085 223.18 45.205 ;
        RECT  215.27 0 217.56 191.34 ;
        RECT  220.89 0 223.18 191.34 ;
        RECT  226.51 39.085 234.42 45.205 ;
        RECT  226.51 0 228.8 191.34 ;
        RECT  232.13 0 234.42 191.34 ;
        RECT  237.75 39.085 245.66 45.205 ;
        RECT  237.75 0 240.04 191.34 ;
        RECT  243.37 0 245.66 191.34 ;
        RECT  248.99 39.085 256.9 45.205 ;
        RECT  248.99 0 251.28 191.34 ;
        RECT  254.61 0 256.9 191.34 ;
        RECT  260.23 39.085 268.14 45.205 ;
        RECT  260.23 0 262.52 191.34 ;
        RECT  265.85 0 268.14 191.34 ;
        RECT  271.47 39.085 279.38 45.205 ;
        RECT  271.47 0 273.76 191.34 ;
        RECT  277.09 0 279.38 191.34 ;
        RECT  282.71 39.085 290.62 45.205 ;
        RECT  282.71 0 285 191.34 ;
        RECT  288.33 0 290.62 191.34 ;
        RECT  293.95 39.085 301.86 45.205 ;
        RECT  293.95 0 296.24 191.34 ;
        RECT  299.57 0 301.86 191.34 ;
        RECT  305.19 39.085 313.1 45.205 ;
        RECT  305.19 0 307.48 191.34 ;
        RECT  310.81 0 313.1 191.34 ;
        RECT  316.43 39.085 324.34 45.205 ;
        RECT  316.43 0 318.72 191.34 ;
        RECT  322.05 0 324.34 191.34 ;
        RECT  327.67 39.085 335.58 45.205 ;
        RECT  327.67 0 329.96 191.34 ;
        RECT  333.29 0 335.58 191.34 ;
        RECT  338.91 39.085 346.82 45.205 ;
        RECT  338.91 0 341.2 191.34 ;
        RECT  344.53 0 346.82 191.34 ;
        RECT  350.15 39.085 358.06 45.205 ;
        RECT  350.15 0 352.44 191.34 ;
        RECT  355.77 0 358.06 191.34 ;
        RECT  361.39 0 372.55 191.34 ;
        RECT  375.88 0 377.7 191.34 ;
        RECT  381.03 0 382.85 191.34 ;
        RECT  386.18 0 388 191.34 ;
        RECT  391.33 0 393.15 191.34 ;
        RECT  396.48 0 398.3 191.34 ;
        RECT  426.42 39.085 434.33 45.205 ;
        RECT  426.42 0 428.71 191.34 ;
        RECT  432.04 0 434.33 191.34 ;
        RECT  437.66 39.085 445.57 45.205 ;
        RECT  437.66 0 439.95 191.34 ;
        RECT  443.28 0 445.57 191.34 ;
        RECT  448.9 39.085 456.81 45.205 ;
        RECT  448.9 0 451.19 191.34 ;
        RECT  454.52 0 456.81 191.34 ;
        RECT  460.14 39.085 468.05 45.205 ;
        RECT  460.14 0 462.43 191.34 ;
        RECT  465.76 0 468.05 191.34 ;
        RECT  471.38 39.085 479.29 45.205 ;
        RECT  471.38 0 473.67 191.34 ;
        RECT  477 0 479.29 191.34 ;
        RECT  482.62 39.085 490.53 45.205 ;
        RECT  482.62 0 484.91 191.34 ;
        RECT  488.24 0 490.53 191.34 ;
        RECT  493.86 39.085 501.77 45.205 ;
        RECT  493.86 0 496.15 191.34 ;
        RECT  499.48 0 501.77 191.34 ;
        RECT  505.1 39.085 513.01 45.205 ;
        RECT  505.1 0 507.39 191.34 ;
        RECT  510.72 0 513.01 191.34 ;
        RECT  516.34 39.085 524.25 45.205 ;
        RECT  516.34 0 518.63 191.34 ;
        RECT  521.96 0 524.25 191.34 ;
        RECT  527.58 39.085 535.49 45.205 ;
        RECT  527.58 0 529.87 191.34 ;
        RECT  533.2 0 535.49 191.34 ;
        RECT  538.82 39.085 546.73 45.205 ;
        RECT  538.82 0 541.11 191.34 ;
        RECT  544.44 0 546.73 191.34 ;
        RECT  550.06 39.085 557.97 45.205 ;
        RECT  550.06 0 552.35 191.34 ;
        RECT  555.68 0 557.97 191.34 ;
        RECT  561.3 39.085 569.21 45.205 ;
        RECT  561.3 0 563.59 191.34 ;
        RECT  566.92 0 569.21 191.34 ;
        RECT  572.54 39.085 580.45 45.205 ;
        RECT  572.54 0 574.83 191.34 ;
        RECT  578.16 0 580.45 191.34 ;
        RECT  583.78 39.085 591.69 45.205 ;
        RECT  583.78 0 586.07 191.34 ;
        RECT  589.4 0 591.69 191.34 ;
        RECT  595.02 39.085 602.93 45.205 ;
        RECT  595.02 0 597.31 191.34 ;
        RECT  600.64 0 602.93 191.34 ;
        RECT  606.26 39.085 614.17 45.205 ;
        RECT  606.26 0 608.55 191.34 ;
        RECT  611.88 0 614.17 191.34 ;
        RECT  617.5 39.085 625.41 45.205 ;
        RECT  617.5 0 619.79 191.34 ;
        RECT  623.12 0 625.41 191.34 ;
        RECT  628.74 39.085 636.65 45.205 ;
        RECT  628.74 0 631.03 191.34 ;
        RECT  634.36 0 636.65 191.34 ;
        RECT  639.98 39.085 647.89 45.205 ;
        RECT  639.98 0 642.27 191.34 ;
        RECT  645.6 0 647.89 191.34 ;
        RECT  651.22 39.085 659.13 45.205 ;
        RECT  651.22 0 653.51 191.34 ;
        RECT  656.84 0 659.13 191.34 ;
        RECT  662.46 39.085 670.37 45.205 ;
        RECT  662.46 0 664.75 191.34 ;
        RECT  668.08 0 670.37 191.34 ;
        RECT  673.7 39.085 681.61 45.205 ;
        RECT  673.7 0 675.99 191.34 ;
        RECT  679.32 0 681.61 191.34 ;
        RECT  684.94 39.085 692.85 45.205 ;
        RECT  684.94 0 687.23 191.34 ;
        RECT  690.56 0 692.85 191.34 ;
        RECT  696.18 39.085 704.09 45.205 ;
        RECT  696.18 0 698.47 191.34 ;
        RECT  701.8 0 704.09 191.34 ;
        RECT  707.42 39.085 715.33 45.205 ;
        RECT  707.42 0 709.71 191.34 ;
        RECT  713.04 0 715.33 191.34 ;
        RECT  718.66 39.085 726.57 45.205 ;
        RECT  718.66 0 720.95 191.34 ;
        RECT  724.28 0 726.57 191.34 ;
        RECT  729.9 39.085 737.81 45.205 ;
        RECT  729.9 0 732.19 191.34 ;
        RECT  735.52 0 737.81 191.34 ;
        RECT  741.14 39.085 749.05 45.205 ;
        RECT  741.14 0 743.43 191.34 ;
        RECT  746.76 0 749.05 191.34 ;
        RECT  752.38 39.085 760.29 45.205 ;
        RECT  752.38 0 754.67 191.34 ;
        RECT  758 0 760.29 191.34 ;
        RECT  763.62 39.085 771.53 45.205 ;
        RECT  763.62 0 765.91 191.34 ;
        RECT  769.24 0 771.53 191.34 ;
        RECT  774.86 39.085 784.48 45.205 ;
        RECT  774.86 0 777.15 191.34 ;
        RECT  780.48 0 784.48 191.34 ;
        RECT  401.63 0 403.45 191.34 ;
        RECT  406.78 0 408.6 191.34 ;
        RECT  411.93 0 423.09 191.34 ;
    END
END RM_IHPSG13_1P_512x64_c2_bm_bist
END LIBRARY
