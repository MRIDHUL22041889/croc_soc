VERSION 5.7 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "|" ;

PROPERTYDEFINITIONS
END PROPERTYDEFINITIONS

SITE sg13g2_ioSite
    CLASS PAD ;
    SYMMETRY R90 ;
    SIZE 1 BY 180 ;
END sg13g2_ioSite

MACRO sg13g2_Corner
    CLASS PAD SPACER ;
    SIZE 180 BY 180 ;
    SYMMETRY X Y R90 ;
    SITE sg13g2_ioSite ;
    PIN iovdd
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal3 ;
              RECT  178 66 180 91.5 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  93.5 178 119 180 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  66 178 91.5 180 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  178 93.5 180 119 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  178 66 180 91.5 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  93.5 178 119 180 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  66 178 91.5 180 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  178 93.5 180 119 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  178 66 180 91.5 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  93.5 178 119 180 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  66 178 91.5 180 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  178 93.5 180 119 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  178 66 180 91.5 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  93.5 178 119 180 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  66 178 91.5 180 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  178 93.5 180 119 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  67.5 178 90 180 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  178 67.5 180 90 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  95 178 117.5 180 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  178 95 180 117.5 ;
        END
    END iovdd
    PIN iovss
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal3 ;
              RECT  178 34.5 180 60 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  7 178 32.5 180 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  178 126 180 134 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  126 178 134 180 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  34.5 178 60 180 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  178 7 180 32.5 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  178 34.5 180 60 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  7 178 32.5 180 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  178 126 180 134 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  126 178 134 180 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  34.5 178 60 180 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  178 7 180 32.5 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  178 34.5 180 60 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  7 178 32.5 180 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  178 126 180 134 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  126 178 134 180 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  34.5 178 60 180 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  178 7 180 32.5 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  178 34.5 180 60 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  7 178 32.5 180 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  178 126 180 134 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  126 178 134 180 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  34.5 178 60 180 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  178 7 180 32.5 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  178 127.5 180 132.5 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  178 36 180 58.5 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  8.5 178 31 180 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  178 8.5 180 31 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  36 178 58.5 180 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  127.5 178 132.5 180 ;
        END
    END iovss
    PIN vdd
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal3 ;
              RECT  160 178.59 178 180 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  178.59 160 180 178 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  178 140 180 155.8 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  140 178 155.8 180 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  178 140 180 158 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  140 178 158 180 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  178 140 180 158 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  140 178 158 180 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal3 ;
              RECT  178 140 180 158 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  140 178 158 180 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  178.59 162.2 180 178 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  162.2 178.59 178 180 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  160 178.59 178 180 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  178.59 160 180 178 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  160 178.59 178 180 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  178.59 160 180 178 ;
        END
    END vss
    OBS
      LAYER Metal1 ;
        RECT  0 0 180 180 ;
      LAYER Metal2 ;
        RECT  0 0 180 180 ;
      LAYER Metal3 ;
        RECT  0 0 180 180 ;
      LAYER Metal4 ;
        RECT  0 0 180 180 ;
      LAYER Metal5 ;
        RECT  0 0 180 180 ;
      LAYER TopMetal1 ;
        RECT  0 0 180 180 ;
      LAYER TopMetal2 ;
        RECT  0 0 180 180 ;
      LAYER Via1 ;
        RECT  0 0 180 180 ;
      LAYER Via2 ;
        RECT  0 0 180 180 ;
    END
END sg13g2_Corner

MACRO sg13g2_Filler200
    CLASS PAD SPACER ;
    SIZE 1 BY 180 ;
    SYMMETRY X Y R90 ;
    SITE sg13g2_ioSite ;
    PIN iovdd
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal3 ;
              RECT  0 66 1 91.5 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  0 93.5 1 119 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 66 1 91.5 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 93.5 1 119 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 66 1 91.5 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 93.5 1 119 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 66 1 91.5 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 93.5 1 119 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 95 1 117.5 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 67.5 1 90 ;
        END
    END iovdd
    PIN iovss
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal3 ;
              RECT  0 7 1 32.5 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  0 126 1 134 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  0 34.5 1 60 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 7 1 32.5 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 126 1 134 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 34.5 1 60 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 7 1 32.5 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 126 1 134 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 34.5 1 60 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 7 1 32.5 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 126 1 134 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 34.5 1 60 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 8.5 1 31 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 127.5 1 132.5 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 36 1 58.5 ;
        END
    END iovss
    PIN vdd
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal3 ;
              RECT  0 160 1 178 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 140 1 155.8 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 140 1 158 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 140 1 158 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal3 ;
              RECT  0 140 1 158 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 162.2 1 178 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 160 1 178 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 160 1 178 ;
        END
    END vss
    OBS
      LAYER Metal1 ;
        RECT  0 0 1 180 ;
      LAYER Metal2 ;
        RECT  0 0 1 180 ;
      LAYER Metal3 ;
        RECT  0 0 80 178 ;
      LAYER Metal4 ;
        RECT  0 0 80 178 ;
      LAYER Metal5 ;
        RECT  0 0 80 178 ;
      LAYER TopMetal1 ;
        RECT  0 0 80 178 ;
      LAYER TopMetal2 ;
        RECT  0 8.5 1 132.5 ;
      LAYER Via1 ;
        RECT  0 0 1 180 ;
      LAYER Via2 ;
        RECT  0 0 1 180 ;
    END
END sg13g2_Filler200

MACRO sg13g2_Filler400
    CLASS PAD SPACER ;
    SIZE 2 BY 180 ;
    SYMMETRY X Y R90 ;
    SITE sg13g2_ioSite ;
    PIN iovdd
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal3 ;
              RECT  0 93.5 2 119 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  0 66 2 91.5 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 93.5 2 119 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 66 2 91.5 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 93.5 2 119 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 66 2 91.5 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 93.5 2 119 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 66 2 91.5 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 67.5 2 90 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 95 2 117.5 ;
        END
    END iovdd
    PIN iovss
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal3 ;
              RECT  0 126 2 134 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  0 7 2 32.5 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  0 34.5 2 60 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 126 2 134 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 7 2 32.5 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 34.5 2 60 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 126 2 134 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 7 2 32.5 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 34.5 2 60 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 126 2 134 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 7 2 32.5 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 34.5 2 60 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 8.5 2 31 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 36 2 58.5 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 127.5 2 132.5 ;
        END
    END iovss
    PIN vdd
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal3 ;
              RECT  0 160 2 178 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 140 2 155.8 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 140 2 158 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 140 2 158 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal3 ;
              RECT  0 140 2 158 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 162.2 2 178 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 160 2 178 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 160 2 178 ;
        END
    END vss
    OBS
      LAYER Metal1 ;
        RECT  0 0 2 180 ;
      LAYER Metal2 ;
        RECT  0 0 2 180 ;
      LAYER Metal3 ;
        RECT  0 0 80 178 ;
      LAYER Metal4 ;
        RECT  0 0 80 178 ;
      LAYER Metal5 ;
        RECT  0 0 80 178 ;
      LAYER TopMetal1 ;
        RECT  0 0 80 178 ;
      LAYER TopMetal2 ;
        RECT  0 8.5 2 132.5 ;
      LAYER Via1 ;
        RECT  0 0 2 180 ;
      LAYER Via2 ;
        RECT  0 0 2 180 ;
    END
END sg13g2_Filler400

MACRO sg13g2_Filler1000
    CLASS PAD SPACER ;
    SIZE 5 BY 180 ;
    SYMMETRY X Y R90 ;
    SITE sg13g2_ioSite ;
    PIN iovdd
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal3 ;
              RECT  0 66 5 91.5 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  0 93.5 5 119 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 66 5 91.5 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 93.5 5 119 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 66 5 91.5 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 93.5 5 119 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 66 5 91.5 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 93.5 5 119 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 95 5 117.5 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 67.5 5 90 ;
        END
    END iovdd
    PIN iovss
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal3 ;
              RECT  0 34.5 5 60 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  0 7 5 32.5 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  0 126 5 134 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 34.5 5 60 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 7 5 32.5 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 126 5 134 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 34.5 5 60 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 7 5 32.5 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 126 5 134 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 34.5 5 60 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 7 5 32.5 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 126 5 134 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 127.5 5 132.5 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 36 5 58.5 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 8.5 5 31 ;
        END
    END iovss
    PIN vdd
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal3 ;
              RECT  0 160 5 178 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 140 5 155.8 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 140 5 158 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 140 5 158 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal3 ;
              RECT  0 140 5 158 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 162.2 5 178 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 160 5 178 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 160 5 178 ;
        END
    END vss
    OBS
      LAYER Metal1 ;
        RECT  0 0 5 180 ;
      LAYER Metal2 ;
        RECT  0 0 5 180 ;
      LAYER Metal3 ;
        RECT  0 0 80 178 ;
      LAYER Metal4 ;
        RECT  0 0 80 178 ;
      LAYER Metal5 ;
        RECT  0 0 80 178 ;
      LAYER TopMetal1 ;
        RECT  0 0 80 178 ;
      LAYER TopMetal2 ;
        RECT  0 8.5 5 132.5 ;
      LAYER Via1 ;
        RECT  0 0 5 180 ;
      LAYER Via2 ;
        RECT  0 0 5 180 ;
    END
END sg13g2_Filler1000

MACRO sg13g2_Filler2000
    CLASS PAD SPACER ;
    SIZE 10 BY 180 ;
    SYMMETRY X Y R90 ;
    SITE sg13g2_ioSite ;
    PIN iovdd
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal3 ;
              RECT  0 66 10 91.5 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  0 93.5 10 119 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 66 10 91.5 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 93.5 10 119 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 66 10 91.5 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 93.5 10 119 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 66 10 91.5 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 93.5 10 119 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 67.5 10 90 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 95 10 117.5 ;
        END
    END iovdd
    PIN iovss
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal3 ;
              RECT  0 126 10 134 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  0 7 10 32.5 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  0 34.5 10 60 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 126 10 134 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 7 10 32.5 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 34.5 10 60 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 126 10 134 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 7 10 32.5 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 34.5 10 60 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 126 10 134 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 7 10 32.5 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 34.5 10 60 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 8.5 10 31 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 36 10 58.5 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 127.5 10 132.5 ;
        END
    END iovss
    PIN vdd
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal3 ;
              RECT  0 160 10 178 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 140 10 155.8 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 140 10 158 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 140 10 158 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal3 ;
              RECT  0 140 10 158 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 162.2 10 178 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 160 10 178 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 160 10 178 ;
        END
    END vss
    OBS
      LAYER Metal1 ;
        RECT  0 0 10 180 ;
      LAYER Metal2 ;
        RECT  0 0 10 180 ;
      LAYER Metal3 ;
        RECT  0 0 80 178 ;
      LAYER Metal4 ;
        RECT  0 0 80 178 ;
      LAYER Metal5 ;
        RECT  0 0 80 178 ;
      LAYER TopMetal1 ;
        RECT  0 0 80 178 ;
      LAYER TopMetal2 ;
        RECT  0 8.5 10 132.5 ;
      LAYER Via1 ;
        RECT  0 0 10 180 ;
      LAYER Via2 ;
        RECT  0 0 10 180 ;
    END
END sg13g2_Filler2000

MACRO sg13g2_Filler4000
    CLASS PAD SPACER ;
    SIZE 20 BY 180 ;
    SYMMETRY X Y R90 ;
    SITE sg13g2_ioSite ;
    PIN iovdd
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal3 ;
              RECT  0 66 20 91.5 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  0 93.5 20 119 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 66 20 91.5 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 93.5 20 119 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 66 20 91.5 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 93.5 20 119 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 66 20 91.5 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 93.5 20 119 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 95 20 117.5 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 67.5 20 90 ;
        END
    END iovdd
    PIN iovss
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal3 ;
              RECT  0 7 20 32.5 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  0 34.5 20 60 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  0 126 20 134 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 7 20 32.5 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 34.5 20 60 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 126 20 134 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 7 20 32.5 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 34.5 20 60 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 126 20 134 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 7 20 32.5 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 34.5 20 60 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 126 20 134 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 127.5 20 132.5 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 36 20 58.5 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 8.5 20 31 ;
        END
    END iovss
    PIN vdd
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal3 ;
              RECT  0 160 20 178 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 140 20 155.8 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 140 20 158 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 140 20 158 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal3 ;
              RECT  0 140 20 158 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 162.2 20 178 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 160 20 178 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 160 20 178 ;
        END
    END vss
    OBS
      LAYER Metal1 ;
        RECT  0 0 20 180 ;
      LAYER Metal2 ;
        RECT  0 0 20 180 ;
      LAYER Metal3 ;
        RECT  0 0 80 178 ;
      LAYER Metal4 ;
        RECT  0 0 80 178 ;
      LAYER Metal5 ;
        RECT  0 0 80 178 ;
      LAYER TopMetal1 ;
        RECT  0 0 80 178 ;
      LAYER TopMetal2 ;
        RECT  0 8.5 20 132.5 ;
      LAYER Via1 ;
        RECT  0 0 20 180 ;
      LAYER Via2 ;
        RECT  0 0 20 180 ;
    END
END sg13g2_Filler4000

MACRO sg13g2_Filler10000
    CLASS PAD SPACER ;
    SIZE 50 BY 180 ;
    SYMMETRY X Y R90 ;
    SITE sg13g2_ioSite ;
    PIN iovdd
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal3 ;
              RECT  0 66 50 91.5 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  0 93.5 50 119 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 66 50 91.5 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 93.5 50 119 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 66 50 91.5 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 93.5 50 119 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 66 50 91.5 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 93.5 50 119 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 95 50 117.5 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 67.5 50 90 ;
        END
    END iovdd
    PIN iovss
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal3 ;
              RECT  0 7 50 32.5 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  0 126 50 134 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  0 34.5 50 60 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 7 50 32.5 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 126 50 134 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 34.5 50 60 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 7 50 32.5 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 126 50 134 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 34.5 50 60 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 7 50 32.5 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 126 50 134 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 34.5 50 60 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 8.5 50 31 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 127.5 50 132.5 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 36 50 58.5 ;
        END
    END iovss
    PIN vdd
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal3 ;
              RECT  0 160 50 178 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 140 50 155.8 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 140 50 158 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 140 50 158 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal3 ;
              RECT  0 140 50 158 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 162.2 50 178 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 160 50 178 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 160 50 178 ;
        END
    END vss
    OBS
      LAYER Metal1 ;
        RECT  0 0 50 180 ;
      LAYER Metal2 ;
        RECT  0 0 50 180 ;
      LAYER Metal3 ;
        RECT  0 0 80 178 ;
      LAYER Metal4 ;
        RECT  0 0 80 178 ;
      LAYER Metal5 ;
        RECT  0 0 80 178 ;
      LAYER TopMetal1 ;
        RECT  0 0 80 178 ;
      LAYER TopMetal2 ;
        RECT  0 8.5 50 132.5 ;
      LAYER Via1 ;
        RECT  0 0 50 180 ;
      LAYER Via2 ;
        RECT  0 0 50 180 ;
    END
END sg13g2_Filler10000

MACRO sg13g2_IOPadIn
    CLASS PAD INPUT ;
    SIZE 80 BY 180 ;
    SYMMETRY X Y R90 ;
    SITE sg13g2_ioSite ;
    PIN iovdd
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal3 ;
              RECT  0 93.5 80 119 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  0 66 80 91.5 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 93.5 80 119 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 66 80 91.5 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 93.5 80 119 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 66 80 91.5 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 93.5 80 119 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 66 80 91.5 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 95 80 117.5 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 67.5 80 90 ;
        END
    END iovdd
    PIN iovss
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal3 ;
              RECT  0 7 80 32.5 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  0 126 80 134 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  0 34.5 80 60 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 7 80 32.5 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 126 80 134 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 34.5 80 60 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 7 80 32.5 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 126 80 134 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 34.5 80 60 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 7 80 32.5 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 126 80 134 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 34.5 80 60 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 36 80 58.5 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 8.5 80 31 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 127.5 80 132.5 ;
        END
    END iovss
    PIN p2c
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal2 ;
              RECT  39.83 157.81 40.12 180 ;
            LAYER Metal3 ;
              RECT  39.725 179.71 40.225 180 ;
        END
    END p2c
    PIN pad
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal2 ;
              RECT  5 0 75 3 ;
            LAYER Metal3 ;
              RECT  5 0 75 3 ;
            LAYER Metal4 ;
              RECT  5 0 75 3 ;
            LAYER Metal5 ;
              RECT  5 0 75 3 ;
            LAYER TopMetal1 ;
              RECT  5 0 75 3 ;
            LAYER TopMetal2 ;
              RECT  5 0 75 3 ;
        END
    END pad
    PIN vdd
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal3 ;
              RECT  0 160 80 178 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 140 80 155.8 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 140 80 158 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 140 80 158 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal3 ;
              RECT  0 140 80 158 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 162.2 80 178 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 160 80 178 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 160 80 178 ;
        END
    END vss
    OBS
      LAYER Metal1 ;
        RECT  0 0 80 180 ;
      LAYER Metal2 ;
        RECT  0 0 80 180 ;
      LAYER Metal3 ;
        RECT  0 0 80 178 ;
      LAYER Metal4 ;
        RECT  0 0 80 178 ;
      LAYER Metal5 ;
        RECT  0 0 80 178 ;
      LAYER TopMetal1 ;
        RECT  0 0 80 178 ;
      LAYER TopMetal2 ;
        RECT  0 0 80 132.5 ;
      LAYER Via1 ;
        RECT  0 0 80 180 ;
      LAYER Via2 ;
        RECT  0 0 80 180 ;
    END
END sg13g2_IOPadIn

MACRO sg13g2_IOPadOut4mA
    CLASS PAD OUTPUT ;
    SIZE 80 BY 180 ;
    SYMMETRY X Y R90 ;
    SITE sg13g2_ioSite ;
    PIN c2p
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal2 ;
              RECT  38.145 167 41.855 180 ;
            LAYER Metal3 ;
              RECT  38.145 179.71 41.855 180 ;
        END
    END c2p
    PIN iovdd
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal3 ;
              RECT  0 93.5 80 119 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  0 66 80 91.5 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 93.5 80 119 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 66 80 91.5 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 93.5 80 119 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 66 80 91.5 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 93.5 80 119 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 66 80 91.5 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 95 80 117.5 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 67.5 80 90 ;
        END
    END iovdd
    PIN iovss
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal3 ;
              RECT  0 7 80 32.5 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  0 126 80 134 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  0 34.5 80 60 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 7 80 32.5 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 126 80 134 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 34.5 80 60 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 7 80 32.5 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 126 80 134 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 34.5 80 60 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 7 80 32.5 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 126 80 134 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 34.5 80 60 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 36 80 58.5 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 8.5 80 31 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 127.5 80 132.5 ;
        END
    END iovss
    PIN pad
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal2 ;
              RECT  5 0 75 3 ;
            LAYER Metal3 ;
              RECT  5 0 75 3 ;
            LAYER Metal4 ;
              RECT  5 0 75 3 ;
            LAYER Metal5 ;
              RECT  5 0 75 3 ;
            LAYER TopMetal1 ;
              RECT  5 0 75 3 ;
            LAYER TopMetal2 ;
              RECT  5 0 75 3 ;
        END
    END pad
    PIN vdd
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal3 ;
              RECT  0 160 80 178 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 140 80 155.8 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 140 80 158 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 140 80 158 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal3 ;
              RECT  0 140 80 158 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 162.2 80 178 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 160 80 178 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 160 80 178 ;
        END
    END vss
    OBS
      LAYER Metal1 ;
        RECT  0 0 80 180 ;
      LAYER Metal2 ;
        RECT  0 0 80 180 ;
      LAYER Metal3 ;
        RECT  0 0 80 178 ;
      LAYER Metal4 ;
        RECT  0 0 80 178 ;
      LAYER Metal5 ;
        RECT  0 0 80 178 ;
      LAYER TopMetal1 ;
        RECT  0 0 80 178 ;
      LAYER TopMetal2 ;
        RECT  0 0 80 132.5 ;
      LAYER Via1 ;
        RECT  0 0 80 180 ;
      LAYER Via2 ;
        RECT  0 0 80 180 ;
    END
END sg13g2_IOPadOut4mA

MACRO sg13g2_IOPadOut16mA
    CLASS PAD OUTPUT ;
    SIZE 80 BY 180 ;
    SYMMETRY X Y R90 ;
    SITE sg13g2_ioSite ;
    PIN c2p
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal2 ;
              RECT  38.145 167 41.855 180 ;
            LAYER Metal3 ;
              RECT  38.145 179.71 41.855 180 ;
        END
    END c2p
    PIN iovdd
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal3 ;
              RECT  0 93.5 80 119 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  0 66 80 91.5 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 93.5 80 119 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 66 80 91.5 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 93.5 80 119 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 66 80 91.5 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 93.5 80 119 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 66 80 91.5 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 95 80 117.5 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 67.5 80 90 ;
        END
    END iovdd
    PIN iovss
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal3 ;
              RECT  0 7 80 32.5 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  0 126 80 134 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  0 34.5 80 60 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 7 80 32.5 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 126 80 134 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 34.5 80 60 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 7 80 32.5 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 126 80 134 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 34.5 80 60 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 7 80 32.5 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 126 80 134 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 34.5 80 60 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 36 80 58.5 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 8.5 80 31 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 127.5 80 132.5 ;
        END
    END iovss
    PIN pad
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal2 ;
              RECT  5 0 75 3 ;
            LAYER Metal3 ;
              RECT  5 0 75 3 ;
            LAYER Metal4 ;
              RECT  5 0 75 3 ;
            LAYER Metal5 ;
              RECT  5 0 75 3 ;
            LAYER TopMetal1 ;
              RECT  5 0 75 3 ;
            LAYER TopMetal2 ;
              RECT  5 0 75 3 ;
        END
    END pad
    PIN vdd
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal3 ;
              RECT  0 160 80 178 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 140 80 155.8 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 140 80 158 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 140 80 158 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal3 ;
              RECT  0 140 80 158 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 162.2 80 178 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 160 80 178 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 160 80 178 ;
        END
    END vss
    OBS
      LAYER Metal1 ;
        RECT  0 0 80 180 ;
      LAYER Metal2 ;
        RECT  0 0 80 180 ;
      LAYER Metal3 ;
        RECT  0 0 80 178 ;
      LAYER Metal4 ;
        RECT  0 0 80 178 ;
      LAYER Metal5 ;
        RECT  0 0 80 178 ;
      LAYER TopMetal1 ;
        RECT  0 0 80 178 ;
      LAYER TopMetal2 ;
        RECT  0 0 80 132.5 ;
      LAYER Via1 ;
        RECT  0 0 80 180 ;
      LAYER Via2 ;
        RECT  0 0 80 180 ;
    END
END sg13g2_IOPadOut16mA

MACRO sg13g2_IOPadOut30mA
    CLASS PAD OUTPUT ;
    SIZE 80 BY 180 ;
    SYMMETRY X Y R90 ;
    SITE sg13g2_ioSite ;
    PIN c2p
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal2 ;
              RECT  38.145 167 41.855 180 ;
            LAYER Metal3 ;
              RECT  38.145 179.71 41.855 180 ;
        END
    END c2p
    PIN iovdd
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal3 ;
              RECT  0 93.5 80 119 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  0 66 80 91.5 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 93.5 80 119 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 66 80 91.5 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 93.5 80 119 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 66 80 91.5 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 93.5 80 119 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 66 80 91.5 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 95 80 117.5 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 67.5 80 90 ;
        END
    END iovdd
    PIN iovss
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal3 ;
              RECT  0 7 80 32.5 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  0 126 80 134 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  0 34.5 80 60 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 7 80 32.5 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 126 80 134 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 34.5 80 60 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 7 80 32.5 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 126 80 134 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 34.5 80 60 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 7 80 32.5 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 126 80 134 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 34.5 80 60 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 36 80 58.5 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 8.5 80 31 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 127.5 80 132.5 ;
        END
    END iovss
    PIN pad
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal2 ;
              RECT  5 0 75 3 ;
            LAYER Metal3 ;
              RECT  5 0 75 3 ;
            LAYER Metal4 ;
              RECT  5 0 75 3 ;
            LAYER Metal5 ;
              RECT  5 0 75 3 ;
            LAYER TopMetal1 ;
              RECT  5 0 75 3 ;
            LAYER TopMetal2 ;
              RECT  5 0 75 3 ;
        END
    END pad
    PIN vdd
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal3 ;
              RECT  0 160 80 178 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 140 80 155.8 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 140 80 158 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 140 80 158 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal3 ;
              RECT  0 140 80 158 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 162.2 80 178 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 160 80 178 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 160 80 178 ;
        END
    END vss
    OBS
      LAYER Metal1 ;
        RECT  0 0 80 180 ;
      LAYER Metal2 ;
        RECT  0 0 80 180 ;
      LAYER Metal3 ;
        RECT  0 0 80 178 ;
      LAYER Metal4 ;
        RECT  0 0 80 178 ;
      LAYER Metal5 ;
        RECT  0 0 80 178 ;
      LAYER TopMetal1 ;
        RECT  0 0 80 178 ;
      LAYER TopMetal2 ;
        RECT  0 0 80 132.5 ;
      LAYER Via1 ;
        RECT  0 0 80 180 ;
      LAYER Via2 ;
        RECT  0 0 80 180 ;
    END
END sg13g2_IOPadOut30mA

MACRO sg13g2_IOPadTriOut4mA
    CLASS PAD OUTPUT ;
    SIZE 80 BY 180 ;
    SYMMETRY X Y R90 ;
    SITE sg13g2_ioSite ;
    PIN c2p
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal2 ;
              RECT  38.33 178.09 38.62 180 ;
            LAYER Metal3 ;
              RECT  38.225 179.71 38.725 180 ;
        END
    END c2p
    PIN c2p_en
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal2 ;
              RECT  41.38 174.045 41.67 180 ;
            LAYER Metal3 ;
              RECT  41.275 179.71 41.775 180 ;
        END
    END c2p_en
    PIN iovdd
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal3 ;
              RECT  0 93.5 80 119 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  0 66 80 91.5 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 93.5 80 119 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 66 80 91.5 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 93.5 80 119 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 66 80 91.5 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 93.5 80 119 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 66 80 91.5 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 95 80 117.5 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 67.5 80 90 ;
        END
    END iovdd
    PIN iovss
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal3 ;
              RECT  0 7 80 32.5 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  0 126 80 134 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  0 34.5 80 60 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 7 80 32.5 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 126 80 134 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 34.5 80 60 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 7 80 32.5 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 126 80 134 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 34.5 80 60 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 7 80 32.5 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 126 80 134 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 34.5 80 60 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 36 80 58.5 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 8.5 80 31 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 127.5 80 132.5 ;
        END
    END iovss
    PIN pad
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal2 ;
              RECT  5 0 75 3 ;
            LAYER Metal3 ;
              RECT  5 0 75 3 ;
            LAYER Metal4 ;
              RECT  5 0 75 3 ;
            LAYER Metal5 ;
              RECT  5 0 75 3 ;
            LAYER TopMetal1 ;
              RECT  5 0 75 3 ;
            LAYER TopMetal2 ;
              RECT  5 0 75 3 ;
        END
    END pad
    PIN vdd
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal3 ;
              RECT  0 160 80 178 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 140 80 155.8 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 140 80 158 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 140 80 158 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal3 ;
              RECT  0 140 80 158 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 162.2 80 178 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 160 80 178 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 160 80 178 ;
        END
    END vss
    OBS
      LAYER Metal1 ;
        RECT  0 0 80 180 ;
      LAYER Metal2 ;
        RECT  0 0 80 180 ;
      LAYER Metal3 ;
        RECT  0 0 80 178 ;
      LAYER Metal4 ;
        RECT  0 0 80 178 ;
      LAYER Metal5 ;
        RECT  0 0 80 178 ;
      LAYER TopMetal1 ;
        RECT  0 0 80 178 ;
      LAYER TopMetal2 ;
        RECT  0 0 80 132.5 ;
      LAYER Via1 ;
        RECT  0 0 80 180 ;
      LAYER Via2 ;
        RECT  0 0 80 180 ;
    END
END sg13g2_IOPadTriOut4mA

MACRO sg13g2_IOPadTriOut16mA
    CLASS PAD OUTPUT ;
    SIZE 80 BY 180 ;
    SYMMETRY X Y R90 ;
    SITE sg13g2_ioSite ;
    PIN c2p
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal2 ;
              RECT  38.33 178.09 38.62 180 ;
            LAYER Metal3 ;
              RECT  38.225 179.71 38.725 180 ;
        END
    END c2p
    PIN c2p_en
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal2 ;
              RECT  41.38 174.045 41.67 180 ;
            LAYER Metal3 ;
              RECT  41.275 179.71 41.775 180 ;
        END
    END c2p_en
    PIN iovdd
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal3 ;
              RECT  0 93.5 80 119 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  0 66 80 91.5 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 93.5 80 119 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 66 80 91.5 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 93.5 80 119 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 66 80 91.5 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 93.5 80 119 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 66 80 91.5 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 95 80 117.5 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 67.5 80 90 ;
        END
    END iovdd
    PIN iovss
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal3 ;
              RECT  0 7 80 32.5 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  0 126 80 134 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  0 34.5 80 60 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 7 80 32.5 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 126 80 134 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 34.5 80 60 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 7 80 32.5 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 126 80 134 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 34.5 80 60 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 7 80 32.5 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 126 80 134 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 34.5 80 60 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 36 80 58.5 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 8.5 80 31 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 127.5 80 132.5 ;
        END
    END iovss
    PIN pad
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal2 ;
              RECT  5 0 75 3 ;
            LAYER Metal3 ;
              RECT  5 0 75 3 ;
            LAYER Metal4 ;
              RECT  5 0 75 3 ;
            LAYER Metal5 ;
              RECT  5 0 75 3 ;
            LAYER TopMetal1 ;
              RECT  5 0 75 3 ;
            LAYER TopMetal2 ;
              RECT  5 0 75 3 ;
        END
    END pad
    PIN vdd
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal3 ;
              RECT  0 160 80 178 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 140 80 155.8 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 140 80 158 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 140 80 158 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal3 ;
              RECT  0 140 80 158 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 162.2 80 178 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 160 80 178 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 160 80 178 ;
        END
    END vss
    OBS
      LAYER Metal1 ;
        RECT  0 0 80 180 ;
      LAYER Metal2 ;
        RECT  0 0 80 180 ;
      LAYER Metal3 ;
        RECT  0 0 80 178 ;
      LAYER Metal4 ;
        RECT  0 0 80 178 ;
      LAYER Metal5 ;
        RECT  0 0 80 178 ;
      LAYER TopMetal1 ;
        RECT  0 0 80 178 ;
      LAYER TopMetal2 ;
        RECT  0 0 80 132.5 ;
      LAYER Via1 ;
        RECT  0 0 80 180 ;
      LAYER Via2 ;
        RECT  0 0 80 180 ;
    END
END sg13g2_IOPadTriOut16mA

MACRO sg13g2_IOPadTriOut30mA
    CLASS PAD OUTPUT ;
    SIZE 80 BY 180 ;
    SYMMETRY X Y R90 ;
    SITE sg13g2_ioSite ;
    PIN c2p
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal2 ;
              RECT  38.33 178.09 38.62 180 ;
            LAYER Metal3 ;
              RECT  38.225 179.71 38.725 180 ;
        END
    END c2p
    PIN c2p_en
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal2 ;
              RECT  41.38 174.045 41.67 180 ;
            LAYER Metal3 ;
              RECT  41.275 179.71 41.775 180 ;
        END
    END c2p_en
    PIN iovdd
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal3 ;
              RECT  0 93.5 80 119 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  0 66 80 91.5 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 93.5 80 119 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 66 80 91.5 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 93.5 80 119 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 66 80 91.5 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 93.5 80 119 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 66 80 91.5 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 95 80 117.5 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 67.5 80 90 ;
        END
    END iovdd
    PIN iovss
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal3 ;
              RECT  0 7 80 32.5 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  0 126 80 134 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  0 34.5 80 60 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 7 80 32.5 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 126 80 134 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 34.5 80 60 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 7 80 32.5 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 126 80 134 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 34.5 80 60 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 7 80 32.5 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 126 80 134 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 34.5 80 60 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 36 80 58.5 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 8.5 80 31 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 127.5 80 132.5 ;
        END
    END iovss
    PIN pad
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal2 ;
              RECT  5 0 75 3 ;
            LAYER Metal3 ;
              RECT  5 0 75 3 ;
            LAYER Metal4 ;
              RECT  5 0 75 3 ;
            LAYER Metal5 ;
              RECT  5 0 75 3 ;
            LAYER TopMetal1 ;
              RECT  5 0 75 3 ;
            LAYER TopMetal2 ;
              RECT  5 0 75 3 ;
        END
    END pad
    PIN vdd
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal3 ;
              RECT  0 160 80 178 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 140 80 155.8 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 140 80 158 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 140 80 158 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal3 ;
              RECT  0 140 80 158 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 162.2 80 178 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 160 80 178 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 160 80 178 ;
        END
    END vss
    OBS
      LAYER Metal1 ;
        RECT  0 0 80 180 ;
      LAYER Metal2 ;
        RECT  0 0 80 180 ;
      LAYER Metal3 ;
        RECT  0 0 80 178 ;
      LAYER Metal4 ;
        RECT  0 0 80 178 ;
      LAYER Metal5 ;
        RECT  0 0 80 178 ;
      LAYER TopMetal1 ;
        RECT  0 0 80 178 ;
      LAYER TopMetal2 ;
        RECT  0 0 80 132.5 ;
      LAYER Via1 ;
        RECT  0 0 80 180 ;
      LAYER Via2 ;
        RECT  0 0 80 180 ;
    END
END sg13g2_IOPadTriOut30mA

MACRO sg13g2_IOPadInOut4mA
    CLASS PAD INOUT ;
    SIZE 80 BY 180 ;
    SYMMETRY X Y R90 ;
    SITE sg13g2_ioSite ;
    PIN c2p
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal2 ;
              RECT  18.33 178.09 18.62 180 ;
            LAYER Metal3 ;
              RECT  18.225 179.71 18.725 180 ;
        END
    END c2p
    PIN c2p_en
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal2 ;
              RECT  21.38 174.045 21.67 180 ;
            LAYER Metal3 ;
              RECT  21.275 179.71 21.775 180 ;
        END
    END c2p_en
    PIN iovdd
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal3 ;
              RECT  0 93.5 80 119 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  0 66 80 91.5 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 93.5 80 119 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 66 80 91.5 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 93.5 80 119 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 66 80 91.5 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 93.5 80 119 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 66 80 91.5 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 95 80 117.5 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 67.5 80 90 ;
        END
    END iovdd
    PIN iovss
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal3 ;
              RECT  0 7 80 32.5 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  0 126 80 134 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  0 34.5 80 60 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 7 80 32.5 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 126 80 134 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 34.5 80 60 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 7 80 32.5 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 126 80 134 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 34.5 80 60 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 7 80 32.5 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 126 80 134 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 34.5 80 60 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 36 80 58.5 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 8.5 80 31 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 127.5 80 132.5 ;
        END
    END iovss
    PIN p2c
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal2 ;
              RECT  59.83 157.81 60.12 180 ;
            LAYER Metal3 ;
              RECT  59.725 179.71 60.225 180 ;
        END
    END p2c
    PIN pad
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal2 ;
              RECT  5 0 75 3 ;
            LAYER Metal3 ;
              RECT  5 0 75 3 ;
            LAYER Metal4 ;
              RECT  5 0 75 3 ;
            LAYER Metal5 ;
              RECT  5 0 75 3 ;
            LAYER TopMetal1 ;
              RECT  5 0 75 3 ;
            LAYER TopMetal2 ;
              RECT  5 0 75 3 ;
        END
    END pad
    PIN vdd
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal3 ;
              RECT  0 160 80 178 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 140 80 155.8 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 140 80 158 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 140 80 158 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal3 ;
              RECT  0 140 80 158 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 162.2 80 178 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 160 80 178 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 160 80 178 ;
        END
    END vss
    OBS
      LAYER Metal1 ;
        RECT  0 0 80 180 ;
      LAYER Metal2 ;
        RECT  0 0 80 180 ;
      LAYER Metal3 ;
        RECT  0 0 80 178 ;
      LAYER Metal4 ;
        RECT  0 0 80 178 ;
      LAYER Metal5 ;
        RECT  0 0 80 178 ;
      LAYER TopMetal1 ;
        RECT  0 0 80 178 ;
      LAYER TopMetal2 ;
        RECT  0 0 80 132.5 ;
      LAYER Via1 ;
        RECT  0 0 80 180 ;
      LAYER Via2 ;
        RECT  0 0 80 180 ;
    END
END sg13g2_IOPadInOut4mA

MACRO sg13g2_IOPadInOut16mA
    CLASS PAD INOUT ;
    SIZE 80 BY 180 ;
    SYMMETRY X Y R90 ;
    SITE sg13g2_ioSite ;
    PIN c2p
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal2 ;
              RECT  18.33 178.09 18.62 180 ;
            LAYER Metal3 ;
              RECT  18.225 179.71 18.725 180 ;
        END
    END c2p
    PIN c2p_en
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal2 ;
              RECT  21.38 174.045 21.67 180 ;
            LAYER Metal3 ;
              RECT  21.275 179.71 21.775 180 ;
        END
    END c2p_en
    PIN iovdd
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal3 ;
              RECT  0 93.5 80 119 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  0 66 80 91.5 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 93.5 80 119 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 66 80 91.5 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 93.5 80 119 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 66 80 91.5 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 93.5 80 119 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 66 80 91.5 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 95 80 117.5 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 67.5 80 90 ;
        END
    END iovdd
    PIN iovss
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal3 ;
              RECT  0 7 80 32.5 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  0 126 80 134 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  0 34.5 80 60 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 7 80 32.5 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 126 80 134 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 34.5 80 60 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 7 80 32.5 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 126 80 134 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 34.5 80 60 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 7 80 32.5 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 126 80 134 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 34.5 80 60 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 36 80 58.5 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 8.5 80 31 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 127.5 80 132.5 ;
        END
    END iovss
    PIN p2c
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal2 ;
              RECT  59.83 157.81 60.12 180 ;
            LAYER Metal3 ;
              RECT  59.725 179.71 60.225 180 ;
        END
    END p2c
    PIN pad
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal2 ;
              RECT  5 0 75 3 ;
            LAYER Metal3 ;
              RECT  5 0 75 3 ;
            LAYER Metal4 ;
              RECT  5 0 75 3 ;
            LAYER Metal5 ;
              RECT  5 0 75 3 ;
            LAYER TopMetal1 ;
              RECT  5 0 75 3 ;
            LAYER TopMetal2 ;
              RECT  5 0 75 3 ;
        END
    END pad
    PIN vdd
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal3 ;
              RECT  0 160 80 178 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 140 80 155.8 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 140 80 158 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 140 80 158 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal3 ;
              RECT  0 140 80 158 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 162.2 80 178 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 160 80 178 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 160 80 178 ;
        END
    END vss
    OBS
      LAYER Metal1 ;
        RECT  0 0 80 180 ;
      LAYER Metal2 ;
        RECT  0 0 80 180 ;
      LAYER Metal3 ;
        RECT  0 0 80 178 ;
      LAYER Metal4 ;
        RECT  0 0 80 178 ;
      LAYER Metal5 ;
        RECT  0 0 80 178 ;
      LAYER TopMetal1 ;
        RECT  0 0 80 178 ;
      LAYER TopMetal2 ;
        RECT  0 0 80 132.5 ;
      LAYER Via1 ;
        RECT  0 0 80 180 ;
      LAYER Via2 ;
        RECT  0 0 80 180 ;
    END
END sg13g2_IOPadInOut16mA

MACRO sg13g2_IOPadInOut30mA
    CLASS PAD INOUT ;
    SIZE 80 BY 180 ;
    SYMMETRY X Y R90 ;
    SITE sg13g2_ioSite ;
    PIN c2p
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal2 ;
              RECT  18.33 178.09 18.62 180 ;
            LAYER Metal3 ;
              RECT  18.225 179.71 18.725 180 ;
        END
    END c2p
    PIN c2p_en
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal2 ;
              RECT  21.38 174.045 21.67 180 ;
            LAYER Metal3 ;
              RECT  21.275 179.71 21.775 180 ;
        END
    END c2p_en
    PIN iovdd
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal3 ;
              RECT  0 93.5 80 119 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  0 66 80 91.5 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 93.5 80 119 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 66 80 91.5 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 93.5 80 119 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 66 80 91.5 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 93.5 80 119 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 66 80 91.5 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 95 80 117.5 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 67.5 80 90 ;
        END
    END iovdd
    PIN iovss
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal3 ;
              RECT  0 7 80 32.5 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  0 126 80 134 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  0 34.5 80 60 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 7 80 32.5 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 126 80 134 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 34.5 80 60 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 7 80 32.5 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 126 80 134 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 34.5 80 60 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 7 80 32.5 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 126 80 134 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 34.5 80 60 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 36 80 58.5 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 8.5 80 31 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 127.5 80 132.5 ;
        END
    END iovss
    PIN p2c
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal2 ;
              RECT  59.83 157.81 60.12 180 ;
            LAYER Metal3 ;
              RECT  59.725 179.71 60.225 180 ;
        END
    END p2c
    PIN pad
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal2 ;
              RECT  5 0 75 3 ;
            LAYER Metal3 ;
              RECT  5 0 75 3 ;
            LAYER Metal4 ;
              RECT  5 0 75 3 ;
            LAYER Metal5 ;
              RECT  5 0 75 3 ;
            LAYER TopMetal1 ;
              RECT  5 0 75 3 ;
            LAYER TopMetal2 ;
              RECT  5 0 75 3 ;
        END
    END pad
    PIN vdd
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal3 ;
              RECT  0 160 80 178 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 140 80 155.8 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 140 80 158 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 140 80 158 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal3 ;
              RECT  0 140 80 158 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 162.2 80 178 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 160 80 178 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 160 80 178 ;
        END
    END vss
    OBS
      LAYER Metal1 ;
        RECT  0 0 80 180 ;
      LAYER Metal2 ;
        RECT  0 0 80 180 ;
      LAYER Metal3 ;
        RECT  0 0 80 178 ;
      LAYER Metal4 ;
        RECT  0 0 80 178 ;
      LAYER Metal5 ;
        RECT  0 0 80 178 ;
      LAYER TopMetal1 ;
        RECT  0 0 80 178 ;
      LAYER TopMetal2 ;
        RECT  0 0 80 132.5 ;
      LAYER Via1 ;
        RECT  0 0 80 180 ;
      LAYER Via2 ;
        RECT  0 0 80 180 ;
    END
END sg13g2_IOPadInOut30mA

MACRO sg13g2_IOPadAnalog
    CLASS PAD INOUT ;
    SIZE 80 BY 180 ;
    SYMMETRY X Y R90 ;
    SITE sg13g2_ioSite ;
    PIN iovdd
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal3 ;
              RECT  0 93.5 80 119 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  0 66 80 91.5 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 93.5 80 119 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 66 80 91.5 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 93.5 80 119 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 66 80 91.5 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 93.5 80 119 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 66 80 91.5 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 95 80 117.5 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 67.5 80 90 ;
        END
    END iovdd
    PIN iovss
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal3 ;
              RECT  0 7 80 32.5 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  0 126 80 134 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  0 34.5 80 60 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 7 80 32.5 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 126 80 134 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 34.5 80 60 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 7 80 32.5 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 126 80 134 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 34.5 80 60 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 7 80 32.5 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 126 80 134 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 34.5 80 60 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 36 80 58.5 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 8.5 80 31 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 127.5 80 132.5 ;
        END
    END iovss
    PIN pad
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal2 ;
              RECT  26.105 179 50.875 180 ;
            LAYER Metal3 ;
              RECT  26.105 179.71 50.875 180 ;
        END
        PORT
            LAYER Metal2 ;
              RECT  5 0 75 3 ;
            LAYER Metal3 ;
              RECT  5 0 75 3 ;
            LAYER Metal4 ;
              RECT  5 0 75 3 ;
            LAYER Metal5 ;
              RECT  5 0 75 3 ;
            LAYER TopMetal1 ;
              RECT  5 0 75 3 ;
            LAYER TopMetal2 ;
              RECT  5 0 75 3 ;
        END
    END pad
    PIN padres
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal2 ;
              RECT  57.46 147.18 57.75 180 ;
            LAYER Metal3 ;
              RECT  57.355 179.71 57.855 180 ;
        END
    END padres
    PIN vdd
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal3 ;
              RECT  0 160 80 178 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 140 80 155.8 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 140 80 158 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 140 80 158 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal3 ;
              RECT  0 140 80 158 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 162.2 80 178 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 160 80 178 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 160 80 178 ;
        END
    END vss
    OBS
      LAYER Metal1 ;
        RECT  0 0 80 180 ;
      LAYER Metal2 ;
        RECT  0 0 80 180 ;
      LAYER Metal3 ;
        RECT  0 0 80 178 ;
      LAYER Metal4 ;
        RECT  0 0 80 178 ;
      LAYER Metal5 ;
        RECT  0 0 80 178 ;
      LAYER TopMetal1 ;
        RECT  0 0 80 178 ;
      LAYER TopMetal2 ;
        RECT  0 0 80 132.5 ;
      LAYER Via1 ;
        RECT  0 0 80 180 ;
      LAYER Via2 ;
        RECT  0 0 80 180 ;
    END
END sg13g2_IOPadAnalog

MACRO sg13g2_IOPadIOVss
    CLASS PAD POWER ;
    SIZE 80 BY 180 ;
    SYMMETRY X Y R90 ;
    SITE sg13g2_ioSite ;
    PIN iovdd
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal3 ;
              RECT  0 93.5 80 119 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  0 66 80 91.5 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 93.5 80 119 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 66 80 91.5 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 93.5 80 119 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 66 80 91.5 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 93.5 80 119 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 66 80 91.5 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 95 80 117.5 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 67.5 80 90 ;
        END
    END iovdd
    PIN iovss
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal2 ;
              RECT  5 0 75 3 ;
            LAYER Metal3 ;
              RECT  5 0 75 3 ;
            LAYER Metal4 ;
              RECT  5 0 75 3 ;
            LAYER Metal5 ;
              RECT  5 0 75 3 ;
            LAYER TopMetal1 ;
              RECT  5 0 75 3 ;
            LAYER TopMetal2 ;
              RECT  5 0 75 3 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  0 7 80 32.5 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  0 126 80 134 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  0 34.5 80 60 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 7 80 32.5 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 126 80 134 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 34.5 80 60 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 7 80 32.5 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 126 80 134 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 34.5 80 60 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 7 80 32.5 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 126 80 134 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 34.5 80 60 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 36 80 58.5 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 8.5 80 31 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 127.5 80 132.5 ;
        END
    END iovss
    PIN vdd
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal3 ;
              RECT  0 160 80 178 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 140 80 155.8 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 140 80 158 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 140 80 158 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal3 ;
              RECT  0 140 80 158 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 162.2 80 178 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 160 80 178 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 160 80 178 ;
        END
    END vss
    OBS
      LAYER Metal1 ;
        RECT  0 0 80 180 ;
      LAYER Metal2 ;
        RECT  0 0 80 180 ;
      LAYER Metal3 ;
        RECT  0 0 80 178 ;
      LAYER Metal4 ;
        RECT  0 0 80 178 ;
      LAYER Metal5 ;
        RECT  0 0 80 178 ;
      LAYER TopMetal1 ;
        RECT  0 0 80 178 ;
      LAYER TopMetal2 ;
        RECT  0 0 80 132.5 ;
      LAYER Via1 ;
        RECT  0 0 80 180 ;
      LAYER Via2 ;
        RECT  0 0 80 180 ;
    END
END sg13g2_IOPadIOVss

MACRO sg13g2_IOPadIOVdd
    CLASS PAD POWER ;
    SIZE 80 BY 180 ;
    SYMMETRY X Y R90 ;
    SITE sg13g2_ioSite ;
    PIN iovdd
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal2 ;
              RECT  5 0 75 3 ;
            LAYER Metal3 ;
              RECT  5 0 75 3 ;
            LAYER Metal4 ;
              RECT  5 0 75 3 ;
            LAYER Metal5 ;
              RECT  5 0 75 3 ;
            LAYER TopMetal1 ;
              RECT  5 0 75 3 ;
            LAYER TopMetal2 ;
              RECT  5 0 75 3 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  0 93.5 80 119 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  0 66 80 91.5 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 93.5 80 119 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 66 80 91.5 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 93.5 80 119 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 66 80 91.5 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 93.5 80 119 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 66 80 91.5 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 95 80 117.5 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 67.5 80 90 ;
        END
    END iovdd
    PIN iovss
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal3 ;
              RECT  0 7 80 32.5 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  0 126 80 134 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  0 34.5 80 60 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 7 80 32.5 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 126 80 134 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 34.5 80 60 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 7 80 32.5 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 126 80 134 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 34.5 80 60 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 7 80 32.5 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 126 80 134 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 34.5 80 60 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 36 3.9 58.5 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 8.5 3.9 31 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  76.1 36 80 58.5 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 127.5 80 132.5 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  76.1 8.5 80 31 ;
        END
    END iovss
    PIN vdd
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal3 ;
              RECT  0 160 80 178 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 140 80 155.8 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 140 80 158 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 140 80 158 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal3 ;
              RECT  0 140 80 158 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 162.2 80 178 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 160 80 178 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 160 80 178 ;
        END
    END vss
    OBS
      LAYER Metal1 ;
        RECT  0 0 80 180 ;
      LAYER Metal2 ;
        RECT  0 0 80 180 ;
      LAYER Metal3 ;
        RECT  0 0 80 178 ;
      LAYER Metal4 ;
        RECT  0 0 80 178 ;
      LAYER Metal5 ;
        RECT  0 0 80 178 ;
      LAYER TopMetal1 ;
        RECT  0 0 80 178 ;
      LAYER TopMetal2 ;
        RECT  0 0 80 132.5 ;
      LAYER Via1 ;
        RECT  0 0 80 180 ;
      LAYER Via2 ;
        RECT  0 0 80 180 ;
    END
END sg13g2_IOPadIOVdd

MACRO sg13g2_IOPadVss
    CLASS PAD POWER ;
    SIZE 80 BY 180 ;
    SYMMETRY X Y R90 ;
    SITE sg13g2_ioSite ;
    PIN iovdd
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal3 ;
              RECT  0 93.5 80 119 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  0 66 80 91.5 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 93.5 80 119 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 66 80 91.5 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 93.5 80 119 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 66 80 91.5 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 93.5 80 119 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 66 80 91.5 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 95 80 117.5 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 67.5 80 90 ;
        END
    END iovdd
    PIN iovss
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal3 ;
              RECT  0 7 80 32.5 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  0 126 80 134 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  0 34.5 80 60 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 7 80 32.5 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 126 80 134 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 34.5 80 60 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 7 80 32.5 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 126 80 134 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 34.5 80 60 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 7 80 32.5 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 126 80 134 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 34.5 80 60 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 36 80 58.5 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 8.5 80 31 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 127.5 80 132.5 ;
        END
    END iovss
    PIN vdd
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal3 ;
              RECT  0 160 80 178 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 140 80 155.8 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 140 80 158 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 140 80 158 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal2 ;
              RECT  5 0 75 3 ;
            LAYER Metal3 ;
              RECT  5 0 75 3 ;
            LAYER Metal4 ;
              RECT  5 0 75 3 ;
            LAYER Metal5 ;
              RECT  5 0 75 3 ;
            LAYER TopMetal1 ;
              RECT  5 0 75 3 ;
            LAYER TopMetal2 ;
              RECT  5 0 75 3 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  0 140 80 158 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 162.2 80 178 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 160 80 178 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 160 80 178 ;
        END
    END vss
    OBS
      LAYER Metal1 ;
        RECT  0 0 80 180 ;
      LAYER Metal2 ;
        RECT  0 0 80 180 ;
      LAYER Metal3 ;
        RECT  0 0 80 178 ;
      LAYER Metal4 ;
        RECT  0 0 80 178 ;
      LAYER Metal5 ;
        RECT  0 0 80 178 ;
      LAYER TopMetal1 ;
        RECT  0 0 80 178 ;
      LAYER TopMetal2 ;
        RECT  0 0 80 132.5 ;
      LAYER Via1 ;
        RECT  0 0 80 180 ;
      LAYER Via2 ;
        RECT  0 0 80 180 ;
    END
END sg13g2_IOPadVss

MACRO sg13g2_IOPadVdd
    CLASS PAD POWER ;
    SIZE 80 BY 180 ;
    SYMMETRY X Y R90 ;
    SITE sg13g2_ioSite ;
    PIN iovdd
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal3 ;
              RECT  0 93.5 80 119 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  0 66 80 91.5 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 93.5 80 119 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 66 80 91.5 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 93.5 80 119 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 66 80 91.5 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 93.5 80 119 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 66 80 91.5 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  76.1 67.5 80 90 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  76.1 95 80 117.5 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 95 3.9 117.5 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 67.5 3.9 90 ;
        END
    END iovdd
    PIN iovss
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal3 ;
              RECT  0 7 80 32.5 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  0 126 80 134 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  0 34.5 80 60 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 7 80 32.5 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 126 80 134 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 34.5 80 60 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 7 80 32.5 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 126 80 134 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 34.5 80 60 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 7 80 32.5 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 126 80 134 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 34.5 80 60 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 36 3.9 58.5 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 8.5 3.9 31 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  76.1 127.5 80 132.5 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  76.1 36 80 58.5 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  76.1 8.5 80 31 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  0 127.5 3.9 132.5 ;
        END
    END iovss
    PIN vdd
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal2 ;
              RECT  5 0 75 3 ;
            LAYER Metal3 ;
              RECT  5 0 75 3 ;
            LAYER Metal4 ;
              RECT  5 0 75 3 ;
            LAYER Metal5 ;
              RECT  5 0 75 3 ;
            LAYER TopMetal1 ;
              RECT  5 0 75 3 ;
            LAYER TopMetal2 ;
              RECT  5 0 75 3 ;
        END
        PORT
            LAYER Metal3 ;
              RECT  0 160 80 178 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 140 80 155.8 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 140 80 158 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 140 80 158 ;
        END
        PORT
            LAYER TopMetal2 ;
              RECT  7.5 141.5 72.5 156.5 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal3 ;
              RECT  0 140 80 158 ;
        END
        PORT
            LAYER Metal4 ;
              RECT  0 162.2 80 178 ;
        END
        PORT
            LAYER Metal5 ;
              RECT  0 160 80 178 ;
        END
        PORT
            LAYER TopMetal1 ;
              RECT  0 160 80 178 ;
        END
    END vss
    OBS
      LAYER Metal1 ;
        RECT  0 0 80 180 ;
      LAYER Metal2 ;
        RECT  0 0 80 180 ;
      LAYER Metal3 ;
        RECT  0 0 80 178 ;
      LAYER Metal4 ;
        RECT  0 0 80 178 ;
      LAYER Metal5 ;
        RECT  0 0 80 178 ;
      LAYER TopMetal1 ;
        RECT  0 0 80 178 ;
      LAYER TopMetal2 ;
        RECT  0 0 80 156.5 ;
      LAYER Via1 ;
        RECT  0 0 80 180 ;
      LAYER Via2 ;
        RECT  0 0 80 180 ;
    END
END sg13g2_IOPadVdd
END LIBRARY
